magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 1 21 1303 203
rect 30 -17 64 21
<< locali >>
rect 975 325 1025 425
rect 1143 325 1193 425
rect 1311 325 1352 483
rect 975 291 1352 325
rect 22 215 89 257
rect 207 215 538 257
rect 607 215 860 257
rect 1284 181 1352 291
rect 191 145 1352 181
rect 191 51 257 145
rect 359 51 425 145
rect 631 51 697 145
rect 799 51 865 145
rect 967 51 1033 145
rect 1135 51 1201 145
rect 1303 63 1352 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 22 325 81 493
rect 115 359 165 527
rect 199 393 249 493
rect 283 427 333 527
rect 367 393 417 493
rect 451 427 501 527
rect 555 459 1277 493
rect 555 427 605 459
rect 723 427 773 459
rect 639 393 689 425
rect 807 393 857 425
rect 199 359 857 393
rect 891 359 941 459
rect 1059 359 1109 459
rect 1227 359 1277 459
rect 22 291 941 325
rect 123 181 157 291
rect 907 257 941 291
rect 907 215 1225 257
rect 22 147 157 181
rect 22 51 89 147
rect 123 17 157 111
rect 291 17 325 111
rect 459 17 597 111
rect 731 17 765 111
rect 899 17 933 111
rect 1067 17 1101 111
rect 1235 17 1269 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< labels >>
rlabel locali s 207 215 538 257 6 A
port 1 nsew signal input
rlabel locali s 607 215 860 257 6 B
port 2 nsew signal input
rlabel locali s 22 215 89 257 6 C_N
port 3 nsew signal input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1303 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1303 63 1352 145 6 Y
port 8 nsew signal output
rlabel locali s 1135 51 1201 145 6 Y
port 8 nsew signal output
rlabel locali s 967 51 1033 145 6 Y
port 8 nsew signal output
rlabel locali s 799 51 865 145 6 Y
port 8 nsew signal output
rlabel locali s 631 51 697 145 6 Y
port 8 nsew signal output
rlabel locali s 359 51 425 145 6 Y
port 8 nsew signal output
rlabel locali s 191 51 257 145 6 Y
port 8 nsew signal output
rlabel locali s 191 145 1352 181 6 Y
port 8 nsew signal output
rlabel locali s 1284 181 1352 291 6 Y
port 8 nsew signal output
rlabel locali s 975 291 1352 325 6 Y
port 8 nsew signal output
rlabel locali s 1311 325 1352 483 6 Y
port 8 nsew signal output
rlabel locali s 1143 325 1193 425 6 Y
port 8 nsew signal output
rlabel locali s 975 325 1025 425 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1380 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1128116
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1118016
<< end >>
