magic
tech sky130A
magscale 1 2
timestamp 1679235063
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_0
timestamp 1679235063
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_5595914180890  sky130_fd_pr__hvdfm1sd2__example_5595914180890_1
timestamp 1679235063
transform 1 0 200 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 31290690
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 31289764
<< end >>
