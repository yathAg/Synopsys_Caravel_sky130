magic
tech sky130A
timestamp 1679235063
<< properties >>
string GDS_END 49572
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 49248
<< end >>
