magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 498 582
<< pwell >>
rect 14 21 396 157
rect 29 -17 63 21
<< locali >>
rect 17 237 86 391
rect 358 367 443 493
rect 188 216 254 323
rect 390 105 443 367
rect 312 51 443 105
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 32 435 86 527
rect 120 427 173 493
rect 120 190 154 427
rect 222 367 324 527
rect 37 182 154 190
rect 290 182 356 287
rect 37 139 356 182
rect 37 56 98 139
rect 190 17 278 105
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
<< metal1 >>
rect 0 561 460 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 460 561
rect 0 496 460 527
rect 0 17 460 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 460 17
rect 0 -48 460 -17
<< labels >>
rlabel locali s 17 237 86 391 6 A
port 1 nsew signal input
rlabel locali s 188 216 254 323 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 460 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 14 21 396 157 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 498 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 460 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 312 51 443 105 6 X
port 7 nsew signal output
rlabel locali s 390 105 443 367 6 X
port 7 nsew signal output
rlabel locali s 358 367 443 493 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 460 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3825412
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3820990
<< end >>
