magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -36 679 294 1471
<< poly >>
rect 114 703 144 937
rect 48 687 144 703
rect 48 653 64 687
rect 98 653 144 687
rect 48 637 144 653
rect 114 329 144 637
<< polycont >>
rect 64 653 98 687
<< locali >>
rect 0 1397 258 1431
rect 62 1130 96 1397
rect 64 687 98 703
rect 64 637 98 653
rect 162 687 196 1196
rect 162 653 213 687
rect 162 144 196 653
rect 62 17 96 144
rect 0 -17 258 17
use contact_12  contact_12_0
timestamp 1679235063
transform 1 0 48 0 1 637
box 0 0 1 1
use nmos_m4_w1_260_sli_dli_da_p  nmos_m4_w1_260_sli_dli_da_p_0
timestamp 1679235063
transform 1 0 54 0 1 51
box -26 -26 176 278
use pmos_m4_w2_000_sli_dli_da_p  pmos_m4_w2_000_sli_dli_da_p_0
timestamp 1679235063
transform 1 0 54 0 1 963
box -59 -54 209 454
<< labels >>
rlabel locali s 196 670 196 670 4 Z
port 2 nsew
rlabel locali s 81 670 81 670 4 A
port 1 nsew
rlabel locali s 129 1414 129 1414 4 vdd
port 3 nsew
rlabel locali s 129 0 129 0 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 258 1414
string GDS_END 4083882
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4082488
<< end >>
