magic
tech sky130A
magscale 1 2
timestamp 1679235063
use sky130_fd_pr__dfl1sd__example_55959141808510  sky130_fd_pr__dfl1sd__example_55959141808510_0
timestamp 1679235063
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808280  sky130_fd_pr__hvdfl1sd__example_55959141808280_0
timestamp 1679235063
transform -1 0 0 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 48471556
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48470632
<< end >>
