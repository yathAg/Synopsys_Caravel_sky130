magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< locali >>
rect 175 1140 182 1174
rect 216 1140 254 1174
rect 288 1140 326 1174
rect 360 1140 398 1174
rect 432 1140 470 1174
rect 504 1140 542 1174
rect 576 1140 581 1174
rect 175 20 182 54
rect 216 20 254 54
rect 288 20 326 54
rect 360 20 398 54
rect 432 20 470 54
rect 504 20 542 54
rect 576 20 581 54
<< viali >>
rect 182 1140 216 1174
rect 254 1140 288 1174
rect 326 1140 360 1174
rect 398 1140 432 1174
rect 470 1140 504 1174
rect 542 1140 576 1174
rect 182 20 216 54
rect 254 20 288 54
rect 326 20 360 54
rect 398 20 432 54
rect 470 20 504 54
rect 542 20 576 54
<< obsli1 >>
rect 38 1010 72 1048
rect 38 938 72 976
rect 38 866 72 904
rect 38 794 72 832
rect 38 722 72 760
rect 38 650 72 688
rect 38 578 72 616
rect 38 506 72 544
rect 38 434 72 472
rect 38 362 72 400
rect 38 290 72 328
rect 38 218 72 256
rect 38 112 72 184
rect 149 88 183 1106
rect 255 88 289 1106
rect 361 88 395 1106
rect 467 88 501 1106
rect 573 88 607 1106
rect 684 1010 718 1048
rect 684 938 718 976
rect 684 866 718 904
rect 684 794 718 832
rect 684 722 718 760
rect 684 650 718 688
rect 684 578 718 616
rect 684 506 718 544
rect 684 434 718 472
rect 684 362 718 400
rect 684 290 718 328
rect 684 218 718 256
rect 684 112 718 184
<< obsli1c >>
rect 38 1048 72 1082
rect 38 976 72 1010
rect 38 904 72 938
rect 38 832 72 866
rect 38 760 72 794
rect 38 688 72 722
rect 38 616 72 650
rect 38 544 72 578
rect 38 472 72 506
rect 38 400 72 434
rect 38 328 72 362
rect 38 256 72 290
rect 38 184 72 218
rect 684 1048 718 1082
rect 684 976 718 1010
rect 684 904 718 938
rect 684 832 718 866
rect 684 760 718 794
rect 684 688 718 722
rect 684 616 718 650
rect 684 544 718 578
rect 684 472 718 506
rect 684 400 718 434
rect 684 328 718 362
rect 684 256 718 290
rect 684 184 718 218
<< metal1 >>
rect 170 1174 588 1194
rect 170 1140 182 1174
rect 216 1140 254 1174
rect 288 1140 326 1174
rect 360 1140 398 1174
rect 432 1140 470 1174
rect 504 1140 542 1174
rect 576 1140 588 1174
rect 170 1128 588 1140
rect 26 1082 84 1094
rect 26 1048 38 1082
rect 72 1048 84 1082
rect 26 1010 84 1048
rect 26 976 38 1010
rect 72 976 84 1010
rect 26 938 84 976
rect 26 904 38 938
rect 72 904 84 938
rect 26 866 84 904
rect 26 832 38 866
rect 72 832 84 866
rect 26 794 84 832
rect 26 760 38 794
rect 72 760 84 794
rect 26 722 84 760
rect 26 688 38 722
rect 72 688 84 722
rect 26 650 84 688
rect 26 616 38 650
rect 72 616 84 650
rect 26 578 84 616
rect 26 544 38 578
rect 72 544 84 578
rect 26 506 84 544
rect 26 472 38 506
rect 72 472 84 506
rect 26 434 84 472
rect 26 400 38 434
rect 72 400 84 434
rect 26 362 84 400
rect 26 328 38 362
rect 72 328 84 362
rect 26 290 84 328
rect 26 256 38 290
rect 72 256 84 290
rect 26 218 84 256
rect 26 184 38 218
rect 72 184 84 218
rect 26 100 84 184
rect 672 1082 730 1094
rect 672 1048 684 1082
rect 718 1048 730 1082
rect 672 1010 730 1048
rect 672 976 684 1010
rect 718 976 730 1010
rect 672 938 730 976
rect 672 904 684 938
rect 718 904 730 938
rect 672 866 730 904
rect 672 832 684 866
rect 718 832 730 866
rect 672 794 730 832
rect 672 760 684 794
rect 718 760 730 794
rect 672 722 730 760
rect 672 688 684 722
rect 718 688 730 722
rect 672 650 730 688
rect 672 616 684 650
rect 718 616 730 650
rect 672 578 730 616
rect 672 544 684 578
rect 718 544 730 578
rect 672 506 730 544
rect 672 472 684 506
rect 718 472 730 506
rect 672 434 730 472
rect 672 400 684 434
rect 718 400 730 434
rect 672 362 730 400
rect 672 328 684 362
rect 718 328 730 362
rect 672 290 730 328
rect 672 256 684 290
rect 718 256 730 290
rect 672 218 730 256
rect 672 184 684 218
rect 718 184 730 218
rect 672 100 730 184
rect 170 54 588 66
rect 170 20 182 54
rect 216 20 254 54
rect 288 20 326 54
rect 360 20 398 54
rect 432 20 470 54
rect 504 20 542 54
rect 576 20 588 54
rect 170 0 588 20
<< obsm1 >>
rect 140 100 192 1094
rect 246 100 298 1094
rect 352 100 404 1094
rect 458 100 510 1094
rect 564 100 616 1094
<< metal2 >>
rect 0 622 756 1094
rect 0 100 756 572
<< labels >>
rlabel metal2 s 0 622 756 1094 6 DRAIN
port 1 nsew
rlabel viali s 542 1140 576 1174 6 GATE
port 2 nsew
rlabel viali s 542 20 576 54 6 GATE
port 2 nsew
rlabel viali s 470 1140 504 1174 6 GATE
port 2 nsew
rlabel viali s 470 20 504 54 6 GATE
port 2 nsew
rlabel viali s 398 1140 432 1174 6 GATE
port 2 nsew
rlabel viali s 398 20 432 54 6 GATE
port 2 nsew
rlabel viali s 326 1140 360 1174 6 GATE
port 2 nsew
rlabel viali s 326 20 360 54 6 GATE
port 2 nsew
rlabel viali s 254 1140 288 1174 6 GATE
port 2 nsew
rlabel viali s 254 20 288 54 6 GATE
port 2 nsew
rlabel viali s 182 1140 216 1174 6 GATE
port 2 nsew
rlabel viali s 182 20 216 54 6 GATE
port 2 nsew
rlabel locali s 175 1140 581 1174 6 GATE
port 2 nsew
rlabel locali s 175 20 581 54 6 GATE
port 2 nsew
rlabel metal1 s 170 1128 588 1194 6 GATE
port 2 nsew
rlabel metal1 s 170 0 588 66 6 GATE
port 2 nsew
rlabel metal2 s 0 100 756 572 6 SOURCE
port 3 nsew
rlabel metal1 s 26 100 84 1094 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 672 100 730 1094 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 756 1194
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5515070
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5492788
<< end >>
