magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< metal1 >>
rect 104 5496 150 5750
rect 1352 5496 1398 5750
rect 2600 5496 2646 5750
rect 3848 5496 3894 5750
rect 5096 5496 5142 5750
rect 6344 5496 6390 5750
rect 7592 5496 7638 5750
rect 8840 5496 8886 5750
rect 10088 5496 10134 5750
rect 11336 5496 11382 5750
rect 12584 5496 12630 5750
rect 13832 5496 13878 5750
rect 15080 5496 15126 5750
rect 16328 5496 16374 5750
rect 17576 5496 17622 5750
rect 18824 5496 18870 5750
rect 20072 5496 20118 5750
rect 21320 5496 21366 5750
rect 22568 5496 22614 5750
rect 23816 5496 23862 5750
rect 25064 5496 25110 5750
rect 26312 5496 26358 5750
rect 27560 5496 27606 5750
rect 28808 5496 28854 5750
rect 30056 5496 30102 5750
rect 31304 5496 31350 5750
rect 32552 5496 32598 5750
rect 33800 5496 33846 5750
rect 35048 5496 35094 5750
rect 36296 5496 36342 5750
rect 37544 5496 37590 5750
rect 38792 5496 38838 5750
rect 199 3428 227 3494
rect 80 3400 227 3428
rect 80 2994 108 3400
rect 272 3348 300 3494
rect 1447 3428 1475 3494
rect 1328 3400 1475 3428
rect 272 3320 572 3348
rect 544 3118 572 3320
rect 1328 2994 1356 3400
rect 1520 3348 1548 3494
rect 2695 3428 2723 3494
rect 2576 3400 2723 3428
rect 1520 3320 1820 3348
rect 1792 3118 1820 3320
rect 2576 2994 2604 3400
rect 2768 3348 2796 3494
rect 3943 3428 3971 3494
rect 3824 3400 3971 3428
rect 2768 3320 3068 3348
rect 3040 3118 3068 3320
rect 3824 2994 3852 3400
rect 4016 3348 4044 3494
rect 5191 3428 5219 3494
rect 5072 3400 5219 3428
rect 4016 3320 4316 3348
rect 4288 3118 4316 3320
rect 5072 2994 5100 3400
rect 5264 3348 5292 3494
rect 6439 3428 6467 3494
rect 6320 3400 6467 3428
rect 5264 3320 5564 3348
rect 5536 3118 5564 3320
rect 6320 2994 6348 3400
rect 6512 3348 6540 3494
rect 7687 3428 7715 3494
rect 7568 3400 7715 3428
rect 6512 3320 6812 3348
rect 6784 3118 6812 3320
rect 7568 2994 7596 3400
rect 7760 3348 7788 3494
rect 8935 3428 8963 3494
rect 8816 3400 8963 3428
rect 7760 3320 8060 3348
rect 8032 3118 8060 3320
rect 8816 2994 8844 3400
rect 9008 3348 9036 3494
rect 10183 3428 10211 3494
rect 10064 3400 10211 3428
rect 9008 3320 9308 3348
rect 9280 3118 9308 3320
rect 10064 2994 10092 3400
rect 10256 3348 10284 3494
rect 11431 3428 11459 3494
rect 11312 3400 11459 3428
rect 10256 3320 10556 3348
rect 10528 3118 10556 3320
rect 11312 2994 11340 3400
rect 11504 3348 11532 3494
rect 12679 3428 12707 3494
rect 12560 3400 12707 3428
rect 11504 3320 11804 3348
rect 11776 3118 11804 3320
rect 12560 2994 12588 3400
rect 12752 3348 12780 3494
rect 13927 3428 13955 3494
rect 13808 3400 13955 3428
rect 12752 3320 13052 3348
rect 13024 3118 13052 3320
rect 13808 2994 13836 3400
rect 14000 3348 14028 3494
rect 15175 3428 15203 3494
rect 15056 3400 15203 3428
rect 14000 3320 14300 3348
rect 14272 3118 14300 3320
rect 15056 2994 15084 3400
rect 15248 3348 15276 3494
rect 16423 3428 16451 3494
rect 16304 3400 16451 3428
rect 15248 3320 15548 3348
rect 15520 3118 15548 3320
rect 16304 2994 16332 3400
rect 16496 3348 16524 3494
rect 17671 3428 17699 3494
rect 17552 3400 17699 3428
rect 16496 3320 16796 3348
rect 16768 3118 16796 3320
rect 17552 2994 17580 3400
rect 17744 3348 17772 3494
rect 18919 3428 18947 3494
rect 18800 3400 18947 3428
rect 17744 3320 18044 3348
rect 18016 3118 18044 3320
rect 18800 2994 18828 3400
rect 18992 3348 19020 3494
rect 20167 3428 20195 3494
rect 20048 3400 20195 3428
rect 18992 3320 19292 3348
rect 19264 3118 19292 3320
rect 20048 2994 20076 3400
rect 20240 3348 20268 3494
rect 21415 3428 21443 3494
rect 21296 3400 21443 3428
rect 20240 3320 20540 3348
rect 20512 3118 20540 3320
rect 21296 2994 21324 3400
rect 21488 3348 21516 3494
rect 22663 3428 22691 3494
rect 22544 3400 22691 3428
rect 21488 3320 21788 3348
rect 21760 3118 21788 3320
rect 22544 2994 22572 3400
rect 22736 3348 22764 3494
rect 23911 3428 23939 3494
rect 23792 3400 23939 3428
rect 22736 3320 23036 3348
rect 23008 3118 23036 3320
rect 23792 2994 23820 3400
rect 23984 3348 24012 3494
rect 25159 3428 25187 3494
rect 25040 3400 25187 3428
rect 23984 3320 24284 3348
rect 24256 3118 24284 3320
rect 25040 2994 25068 3400
rect 25232 3348 25260 3494
rect 26407 3428 26435 3494
rect 26288 3400 26435 3428
rect 25232 3320 25532 3348
rect 25504 3118 25532 3320
rect 26288 2994 26316 3400
rect 26480 3348 26508 3494
rect 27655 3428 27683 3494
rect 27536 3400 27683 3428
rect 26480 3320 26780 3348
rect 26752 3118 26780 3320
rect 27536 2994 27564 3400
rect 27728 3348 27756 3494
rect 28903 3428 28931 3494
rect 28784 3400 28931 3428
rect 27728 3320 28028 3348
rect 28000 3118 28028 3320
rect 28784 2994 28812 3400
rect 28976 3348 29004 3494
rect 30151 3428 30179 3494
rect 30032 3400 30179 3428
rect 28976 3320 29276 3348
rect 29248 3118 29276 3320
rect 30032 2994 30060 3400
rect 30224 3348 30252 3494
rect 31399 3428 31427 3494
rect 31280 3400 31427 3428
rect 30224 3320 30524 3348
rect 30496 3118 30524 3320
rect 31280 2994 31308 3400
rect 31472 3348 31500 3494
rect 32647 3428 32675 3494
rect 32528 3400 32675 3428
rect 31472 3320 31772 3348
rect 31744 3118 31772 3320
rect 32528 2994 32556 3400
rect 32720 3348 32748 3494
rect 33895 3428 33923 3494
rect 33776 3400 33923 3428
rect 32720 3320 33020 3348
rect 32992 3118 33020 3320
rect 33776 2994 33804 3400
rect 33968 3348 33996 3494
rect 35143 3428 35171 3494
rect 35024 3400 35171 3428
rect 33968 3320 34268 3348
rect 34240 3118 34268 3320
rect 35024 2994 35052 3400
rect 35216 3348 35244 3494
rect 36391 3428 36419 3494
rect 36272 3400 36419 3428
rect 35216 3320 35516 3348
rect 35488 3118 35516 3320
rect 36272 2994 36300 3400
rect 36464 3348 36492 3494
rect 37639 3428 37667 3494
rect 37520 3400 37667 3428
rect 36464 3320 36764 3348
rect 36736 3118 36764 3320
rect 37520 2994 37548 3400
rect 37712 3348 37740 3494
rect 38887 3428 38915 3494
rect 38768 3400 38915 3428
rect 37712 3320 38012 3348
rect 37984 3118 38012 3320
rect 38768 2994 38796 3400
rect 38960 3348 38988 3494
rect 38960 3320 39260 3348
rect 39232 3118 39260 3320
rect 80 1192 108 1258
rect 66 1164 108 1192
rect 66 252 94 1164
rect 544 1112 572 1258
rect 530 1084 572 1112
rect 676 1112 704 1258
rect 1140 1192 1168 1258
rect 1328 1192 1356 1258
rect 1140 1164 1182 1192
rect 676 1084 718 1112
rect 530 252 558 1084
rect 690 252 718 1084
rect 1154 252 1182 1164
rect 1314 1164 1356 1192
rect 1314 252 1342 1164
rect 1792 1112 1820 1258
rect 1778 1084 1820 1112
rect 1924 1112 1952 1258
rect 2388 1192 2416 1258
rect 2576 1192 2604 1258
rect 2388 1164 2430 1192
rect 1924 1084 1966 1112
rect 1778 252 1806 1084
rect 1938 252 1966 1084
rect 2402 252 2430 1164
rect 2562 1164 2604 1192
rect 2562 252 2590 1164
rect 3040 1112 3068 1258
rect 3026 1084 3068 1112
rect 3172 1112 3200 1258
rect 3636 1192 3664 1258
rect 3824 1192 3852 1258
rect 3636 1164 3678 1192
rect 3172 1084 3214 1112
rect 3026 252 3054 1084
rect 3186 252 3214 1084
rect 3650 252 3678 1164
rect 3810 1164 3852 1192
rect 3810 252 3838 1164
rect 4288 1112 4316 1258
rect 4274 1084 4316 1112
rect 4420 1112 4448 1258
rect 4884 1192 4912 1258
rect 5072 1192 5100 1258
rect 4884 1164 4926 1192
rect 4420 1084 4462 1112
rect 4274 252 4302 1084
rect 4434 252 4462 1084
rect 4898 252 4926 1164
rect 5058 1164 5100 1192
rect 5058 252 5086 1164
rect 5536 1112 5564 1258
rect 5522 1084 5564 1112
rect 5668 1112 5696 1258
rect 6132 1192 6160 1258
rect 6320 1192 6348 1258
rect 6132 1164 6174 1192
rect 5668 1084 5710 1112
rect 5522 252 5550 1084
rect 5682 252 5710 1084
rect 6146 252 6174 1164
rect 6306 1164 6348 1192
rect 6306 252 6334 1164
rect 6784 1112 6812 1258
rect 6770 1084 6812 1112
rect 6916 1112 6944 1258
rect 7380 1192 7408 1258
rect 7568 1192 7596 1258
rect 7380 1164 7422 1192
rect 6916 1084 6958 1112
rect 6770 252 6798 1084
rect 6930 252 6958 1084
rect 7394 252 7422 1164
rect 7554 1164 7596 1192
rect 7554 252 7582 1164
rect 8032 1112 8060 1258
rect 8018 1084 8060 1112
rect 8164 1112 8192 1258
rect 8628 1192 8656 1258
rect 8816 1192 8844 1258
rect 8628 1164 8670 1192
rect 8164 1084 8206 1112
rect 8018 252 8046 1084
rect 8178 252 8206 1084
rect 8642 252 8670 1164
rect 8802 1164 8844 1192
rect 8802 252 8830 1164
rect 9280 1112 9308 1258
rect 9266 1084 9308 1112
rect 9412 1112 9440 1258
rect 9876 1192 9904 1258
rect 10064 1192 10092 1258
rect 9876 1164 9918 1192
rect 9412 1084 9454 1112
rect 9266 252 9294 1084
rect 9426 252 9454 1084
rect 9890 252 9918 1164
rect 10050 1164 10092 1192
rect 10050 252 10078 1164
rect 10528 1112 10556 1258
rect 10514 1084 10556 1112
rect 10660 1112 10688 1258
rect 11124 1192 11152 1258
rect 11312 1192 11340 1258
rect 11124 1164 11166 1192
rect 10660 1084 10702 1112
rect 10514 252 10542 1084
rect 10674 252 10702 1084
rect 11138 252 11166 1164
rect 11298 1164 11340 1192
rect 11298 252 11326 1164
rect 11776 1112 11804 1258
rect 11762 1084 11804 1112
rect 11908 1112 11936 1258
rect 12372 1192 12400 1258
rect 12560 1192 12588 1258
rect 12372 1164 12414 1192
rect 11908 1084 11950 1112
rect 11762 252 11790 1084
rect 11922 252 11950 1084
rect 12386 252 12414 1164
rect 12546 1164 12588 1192
rect 12546 252 12574 1164
rect 13024 1112 13052 1258
rect 13010 1084 13052 1112
rect 13156 1112 13184 1258
rect 13620 1192 13648 1258
rect 13808 1192 13836 1258
rect 13620 1164 13662 1192
rect 13156 1084 13198 1112
rect 13010 252 13038 1084
rect 13170 252 13198 1084
rect 13634 252 13662 1164
rect 13794 1164 13836 1192
rect 13794 252 13822 1164
rect 14272 1112 14300 1258
rect 14258 1084 14300 1112
rect 14404 1112 14432 1258
rect 14868 1192 14896 1258
rect 15056 1192 15084 1258
rect 14868 1164 14910 1192
rect 14404 1084 14446 1112
rect 14258 252 14286 1084
rect 14418 252 14446 1084
rect 14882 252 14910 1164
rect 15042 1164 15084 1192
rect 15042 252 15070 1164
rect 15520 1112 15548 1258
rect 15506 1084 15548 1112
rect 15652 1112 15680 1258
rect 16116 1192 16144 1258
rect 16304 1192 16332 1258
rect 16116 1164 16158 1192
rect 15652 1084 15694 1112
rect 15506 252 15534 1084
rect 15666 252 15694 1084
rect 16130 252 16158 1164
rect 16290 1164 16332 1192
rect 16290 252 16318 1164
rect 16768 1112 16796 1258
rect 16754 1084 16796 1112
rect 16900 1112 16928 1258
rect 17364 1192 17392 1258
rect 17552 1192 17580 1258
rect 17364 1164 17406 1192
rect 16900 1084 16942 1112
rect 16754 252 16782 1084
rect 16914 252 16942 1084
rect 17378 252 17406 1164
rect 17538 1164 17580 1192
rect 17538 252 17566 1164
rect 18016 1112 18044 1258
rect 18002 1084 18044 1112
rect 18148 1112 18176 1258
rect 18612 1192 18640 1258
rect 18800 1192 18828 1258
rect 18612 1164 18654 1192
rect 18148 1084 18190 1112
rect 18002 252 18030 1084
rect 18162 252 18190 1084
rect 18626 252 18654 1164
rect 18786 1164 18828 1192
rect 18786 252 18814 1164
rect 19264 1112 19292 1258
rect 19250 1084 19292 1112
rect 19396 1112 19424 1258
rect 19860 1192 19888 1258
rect 20048 1192 20076 1258
rect 19860 1164 19902 1192
rect 19396 1084 19438 1112
rect 19250 252 19278 1084
rect 19410 252 19438 1084
rect 19874 252 19902 1164
rect 20034 1164 20076 1192
rect 20034 252 20062 1164
rect 20512 1112 20540 1258
rect 20498 1084 20540 1112
rect 20644 1112 20672 1258
rect 21108 1192 21136 1258
rect 21296 1192 21324 1258
rect 21108 1164 21150 1192
rect 20644 1084 20686 1112
rect 20498 252 20526 1084
rect 20658 252 20686 1084
rect 21122 252 21150 1164
rect 21282 1164 21324 1192
rect 21282 252 21310 1164
rect 21760 1112 21788 1258
rect 21746 1084 21788 1112
rect 21892 1112 21920 1258
rect 22356 1192 22384 1258
rect 22544 1192 22572 1258
rect 22356 1164 22398 1192
rect 21892 1084 21934 1112
rect 21746 252 21774 1084
rect 21906 252 21934 1084
rect 22370 252 22398 1164
rect 22530 1164 22572 1192
rect 22530 252 22558 1164
rect 23008 1112 23036 1258
rect 22994 1084 23036 1112
rect 23140 1112 23168 1258
rect 23604 1192 23632 1258
rect 23792 1192 23820 1258
rect 23604 1164 23646 1192
rect 23140 1084 23182 1112
rect 22994 252 23022 1084
rect 23154 252 23182 1084
rect 23618 252 23646 1164
rect 23778 1164 23820 1192
rect 23778 252 23806 1164
rect 24256 1112 24284 1258
rect 24242 1084 24284 1112
rect 24388 1112 24416 1258
rect 24852 1192 24880 1258
rect 25040 1192 25068 1258
rect 24852 1164 24894 1192
rect 24388 1084 24430 1112
rect 24242 252 24270 1084
rect 24402 252 24430 1084
rect 24866 252 24894 1164
rect 25026 1164 25068 1192
rect 25026 252 25054 1164
rect 25504 1112 25532 1258
rect 25490 1084 25532 1112
rect 25636 1112 25664 1258
rect 26100 1192 26128 1258
rect 26288 1192 26316 1258
rect 26100 1164 26142 1192
rect 25636 1084 25678 1112
rect 25490 252 25518 1084
rect 25650 252 25678 1084
rect 26114 252 26142 1164
rect 26274 1164 26316 1192
rect 26274 252 26302 1164
rect 26752 1112 26780 1258
rect 26738 1084 26780 1112
rect 26884 1112 26912 1258
rect 27348 1192 27376 1258
rect 27536 1192 27564 1258
rect 27348 1164 27390 1192
rect 26884 1084 26926 1112
rect 26738 252 26766 1084
rect 26898 252 26926 1084
rect 27362 252 27390 1164
rect 27522 1164 27564 1192
rect 27522 252 27550 1164
rect 28000 1112 28028 1258
rect 27986 1084 28028 1112
rect 28132 1112 28160 1258
rect 28596 1192 28624 1258
rect 28784 1192 28812 1258
rect 28596 1164 28638 1192
rect 28132 1084 28174 1112
rect 27986 252 28014 1084
rect 28146 252 28174 1084
rect 28610 252 28638 1164
rect 28770 1164 28812 1192
rect 28770 252 28798 1164
rect 29248 1112 29276 1258
rect 29234 1084 29276 1112
rect 29380 1112 29408 1258
rect 29844 1192 29872 1258
rect 30032 1192 30060 1258
rect 29844 1164 29886 1192
rect 29380 1084 29422 1112
rect 29234 252 29262 1084
rect 29394 252 29422 1084
rect 29858 252 29886 1164
rect 30018 1164 30060 1192
rect 30018 252 30046 1164
rect 30496 1112 30524 1258
rect 30482 1084 30524 1112
rect 30628 1112 30656 1258
rect 31092 1192 31120 1258
rect 31280 1192 31308 1258
rect 31092 1164 31134 1192
rect 30628 1084 30670 1112
rect 30482 252 30510 1084
rect 30642 252 30670 1084
rect 31106 252 31134 1164
rect 31266 1164 31308 1192
rect 31266 252 31294 1164
rect 31744 1112 31772 1258
rect 31730 1084 31772 1112
rect 31876 1112 31904 1258
rect 32340 1192 32368 1258
rect 32528 1192 32556 1258
rect 32340 1164 32382 1192
rect 31876 1084 31918 1112
rect 31730 252 31758 1084
rect 31890 252 31918 1084
rect 32354 252 32382 1164
rect 32514 1164 32556 1192
rect 32514 252 32542 1164
rect 32992 1112 33020 1258
rect 32978 1084 33020 1112
rect 33124 1112 33152 1258
rect 33588 1192 33616 1258
rect 33776 1192 33804 1258
rect 33588 1164 33630 1192
rect 33124 1084 33166 1112
rect 32978 252 33006 1084
rect 33138 252 33166 1084
rect 33602 252 33630 1164
rect 33762 1164 33804 1192
rect 33762 252 33790 1164
rect 34240 1112 34268 1258
rect 34226 1084 34268 1112
rect 34372 1112 34400 1258
rect 34836 1192 34864 1258
rect 35024 1192 35052 1258
rect 34836 1164 34878 1192
rect 34372 1084 34414 1112
rect 34226 252 34254 1084
rect 34386 252 34414 1084
rect 34850 252 34878 1164
rect 35010 1164 35052 1192
rect 35010 252 35038 1164
rect 35488 1112 35516 1258
rect 35474 1084 35516 1112
rect 35620 1112 35648 1258
rect 36084 1192 36112 1258
rect 36272 1192 36300 1258
rect 36084 1164 36126 1192
rect 35620 1084 35662 1112
rect 35474 252 35502 1084
rect 35634 252 35662 1084
rect 36098 252 36126 1164
rect 36258 1164 36300 1192
rect 36258 252 36286 1164
rect 36736 1112 36764 1258
rect 36722 1084 36764 1112
rect 36868 1112 36896 1258
rect 37332 1192 37360 1258
rect 37520 1192 37548 1258
rect 37332 1164 37374 1192
rect 36868 1084 36910 1112
rect 36722 252 36750 1084
rect 36882 252 36910 1084
rect 37346 252 37374 1164
rect 37506 1164 37548 1192
rect 37506 252 37534 1164
rect 37984 1112 38012 1258
rect 37970 1084 38012 1112
rect 38116 1112 38144 1258
rect 38580 1192 38608 1258
rect 38768 1192 38796 1258
rect 38580 1164 38622 1192
rect 38116 1084 38158 1112
rect 37970 252 37998 1084
rect 38130 252 38158 1084
rect 38594 252 38622 1164
rect 38754 1164 38796 1192
rect 38754 252 38782 1164
rect 39232 1112 39260 1258
rect 39218 1084 39260 1112
rect 39364 1112 39392 1258
rect 39828 1192 39856 1258
rect 39828 1164 39870 1192
rect 39364 1084 39406 1112
rect 39218 252 39246 1084
rect 39378 252 39406 1084
rect 39842 252 39870 1164
rect 40002 252 40030 1006
rect 40466 252 40494 1006
<< metal3 >>
rect 332 5593 430 5691
rect 1580 5593 1678 5691
rect 2828 5593 2926 5691
rect 4076 5593 4174 5691
rect 5324 5593 5422 5691
rect 6572 5593 6670 5691
rect 7820 5593 7918 5691
rect 9068 5593 9166 5691
rect 10316 5593 10414 5691
rect 11564 5593 11662 5691
rect 12812 5593 12910 5691
rect 14060 5593 14158 5691
rect 15308 5593 15406 5691
rect 16556 5593 16654 5691
rect 17804 5593 17902 5691
rect 19052 5593 19150 5691
rect 20300 5593 20398 5691
rect 21548 5593 21646 5691
rect 22796 5593 22894 5691
rect 24044 5593 24142 5691
rect 25292 5593 25390 5691
rect 26540 5593 26638 5691
rect 27788 5593 27886 5691
rect 29036 5593 29134 5691
rect 30284 5593 30382 5691
rect 31532 5593 31630 5691
rect 32780 5593 32878 5691
rect 34028 5593 34126 5691
rect 35276 5593 35374 5691
rect 36524 5593 36622 5691
rect 37772 5593 37870 5691
rect 39020 5593 39118 5691
rect 332 5271 430 5369
rect 1580 5271 1678 5369
rect 2828 5271 2926 5369
rect 4076 5271 4174 5369
rect 5324 5271 5422 5369
rect 6572 5271 6670 5369
rect 7820 5271 7918 5369
rect 9068 5271 9166 5369
rect 10316 5271 10414 5369
rect 11564 5271 11662 5369
rect 12812 5271 12910 5369
rect 14060 5271 14158 5369
rect 15308 5271 15406 5369
rect 16556 5271 16654 5369
rect 17804 5271 17902 5369
rect 19052 5271 19150 5369
rect 20300 5271 20398 5369
rect 21548 5271 21646 5369
rect 22796 5271 22894 5369
rect 24044 5271 24142 5369
rect 25292 5271 25390 5369
rect 26540 5271 26638 5369
rect 27788 5271 27886 5369
rect 29036 5271 29134 5369
rect 30284 5271 30382 5369
rect 31532 5271 31630 5369
rect 32780 5271 32878 5369
rect 34028 5271 34126 5369
rect 35276 5271 35374 5369
rect 36524 5271 36622 5369
rect 37772 5271 37870 5369
rect 39020 5271 39118 5369
rect 320 4433 418 4531
rect 1568 4433 1666 4531
rect 2816 4433 2914 4531
rect 4064 4433 4162 4531
rect 5312 4433 5410 4531
rect 6560 4433 6658 4531
rect 7808 4433 7906 4531
rect 9056 4433 9154 4531
rect 10304 4433 10402 4531
rect 11552 4433 11650 4531
rect 12800 4433 12898 4531
rect 14048 4433 14146 4531
rect 15296 4433 15394 4531
rect 16544 4433 16642 4531
rect 17792 4433 17890 4531
rect 19040 4433 19138 4531
rect 20288 4433 20386 4531
rect 21536 4433 21634 4531
rect 22784 4433 22882 4531
rect 24032 4433 24130 4531
rect 25280 4433 25378 4531
rect 26528 4433 26626 4531
rect 27776 4433 27874 4531
rect 29024 4433 29122 4531
rect 30272 4433 30370 4531
rect 31520 4433 31618 4531
rect 32768 4433 32866 4531
rect 34016 4433 34114 4531
rect 35264 4433 35362 4531
rect 36512 4433 36610 4531
rect 37760 4433 37858 4531
rect 39008 4433 39106 4531
rect 402 3659 500 3757
rect 1650 3659 1748 3757
rect 2898 3659 2996 3757
rect 4146 3659 4244 3757
rect 5394 3659 5492 3757
rect 6642 3659 6740 3757
rect 7890 3659 7988 3757
rect 9138 3659 9236 3757
rect 10386 3659 10484 3757
rect 11634 3659 11732 3757
rect 12882 3659 12980 3757
rect 14130 3659 14228 3757
rect 15378 3659 15476 3757
rect 16626 3659 16724 3757
rect 17874 3659 17972 3757
rect 19122 3659 19220 3757
rect 20370 3659 20468 3757
rect 21618 3659 21716 3757
rect 22866 3659 22964 3757
rect 24114 3659 24212 3757
rect 25362 3659 25460 3757
rect 26610 3659 26708 3757
rect 27858 3659 27956 3757
rect 29106 3659 29204 3757
rect 30354 3659 30452 3757
rect 31602 3659 31700 3757
rect 32850 3659 32948 3757
rect 34098 3659 34196 3757
rect 35346 3659 35444 3757
rect 36594 3659 36692 3757
rect 37842 3659 37940 3757
rect 39090 3659 39188 3757
rect 0 3526 39936 3586
rect 0 2810 39936 2870
rect 0 2686 39936 2746
rect 575 1886 673 1984
rect 1823 1886 1921 1984
rect 3071 1886 3169 1984
rect 4319 1886 4417 1984
rect 5567 1886 5665 1984
rect 6815 1886 6913 1984
rect 8063 1886 8161 1984
rect 9311 1886 9409 1984
rect 10559 1886 10657 1984
rect 11807 1886 11905 1984
rect 13055 1886 13153 1984
rect 14303 1886 14401 1984
rect 15551 1886 15649 1984
rect 16799 1886 16897 1984
rect 18047 1886 18145 1984
rect 19295 1886 19393 1984
rect 20543 1886 20641 1984
rect 21791 1886 21889 1984
rect 23039 1886 23137 1984
rect 24287 1886 24385 1984
rect 25535 1886 25633 1984
rect 26783 1886 26881 1984
rect 28031 1886 28129 1984
rect 29279 1886 29377 1984
rect 30527 1886 30625 1984
rect 31775 1886 31873 1984
rect 33023 1886 33121 1984
rect 34271 1886 34369 1984
rect 35519 1886 35617 1984
rect 36767 1886 36865 1984
rect 38015 1886 38113 1984
rect 39263 1886 39361 1984
rect 0 951 40560 1011
rect 144 313 242 411
rect 1006 313 1104 411
rect 1392 313 1490 411
rect 2254 313 2352 411
rect 2640 313 2738 411
rect 3502 313 3600 411
rect 3888 313 3986 411
rect 4750 313 4848 411
rect 5136 313 5234 411
rect 5998 313 6096 411
rect 6384 313 6482 411
rect 7246 313 7344 411
rect 7632 313 7730 411
rect 8494 313 8592 411
rect 8880 313 8978 411
rect 9742 313 9840 411
rect 10128 313 10226 411
rect 10990 313 11088 411
rect 11376 313 11474 411
rect 12238 313 12336 411
rect 12624 313 12722 411
rect 13486 313 13584 411
rect 13872 313 13970 411
rect 14734 313 14832 411
rect 15120 313 15218 411
rect 15982 313 16080 411
rect 16368 313 16466 411
rect 17230 313 17328 411
rect 17616 313 17714 411
rect 18478 313 18576 411
rect 18864 313 18962 411
rect 19726 313 19824 411
rect 20112 313 20210 411
rect 20974 313 21072 411
rect 21360 313 21458 411
rect 22222 313 22320 411
rect 22608 313 22706 411
rect 23470 313 23568 411
rect 23856 313 23954 411
rect 24718 313 24816 411
rect 25104 313 25202 411
rect 25966 313 26064 411
rect 26352 313 26450 411
rect 27214 313 27312 411
rect 27600 313 27698 411
rect 28462 313 28560 411
rect 28848 313 28946 411
rect 29710 313 29808 411
rect 30096 313 30194 411
rect 30958 313 31056 411
rect 31344 313 31442 411
rect 32206 313 32304 411
rect 32592 313 32690 411
rect 33454 313 33552 411
rect 33840 313 33938 411
rect 34702 313 34800 411
rect 35088 313 35186 411
rect 35950 313 36048 411
rect 36336 313 36434 411
rect 37198 313 37296 411
rect 37584 313 37682 411
rect 38446 313 38544 411
rect 38832 313 38930 411
rect 39694 313 39792 411
rect 40080 313 40178 411
use precharge_array_0  precharge_array_0_0
timestamp 1679235063
transform 1 0 0 0 -1 1006
box 0 -12 40560 768
use sense_amp_array  sense_amp_array_0
timestamp 1679235063
transform 1 0 0 0 -1 5750
box -160 0 39936 2256
use single_level_column_mux_array_0  single_level_column_mux_array_0_0
timestamp 1679235063
transform 1 0 0 0 -1 3242
box 0 87 39936 1984
<< labels >>
rlabel metal1 s 28831 5623 28831 5623 4 dout_23
port 26 nsew
rlabel metal1 s 26335 5623 26335 5623 4 dout_21
port 24 nsew
rlabel metal1 s 31327 5623 31327 5623 4 dout_25
port 28 nsew
rlabel metal1 s 37567 5623 37567 5623 4 dout_30
port 33 nsew
rlabel metal1 s 23839 5623 23839 5623 4 dout_19
port 22 nsew
rlabel metal1 s 38815 5623 38815 5623 4 dout_31
port 34 nsew
rlabel metal1 s 25087 5623 25087 5623 4 dout_20
port 23 nsew
rlabel metal1 s 35071 5623 35071 5623 4 dout_28
port 31 nsew
rlabel metal1 s 32575 5623 32575 5623 4 dout_26
port 29 nsew
rlabel metal1 s 22591 5623 22591 5623 4 dout_18
port 21 nsew
rlabel metal1 s 27583 5623 27583 5623 4 dout_22
port 25 nsew
rlabel metal1 s 30079 5623 30079 5623 4 dout_24
port 27 nsew
rlabel metal1 s 33823 5623 33823 5623 4 dout_27
port 30 nsew
rlabel metal1 s 36319 5623 36319 5623 4 dout_29
port 32 nsew
rlabel metal1 s 21343 5623 21343 5623 4 dout_17
port 20 nsew
rlabel metal1 s 15103 5623 15103 5623 4 dout_12
port 15 nsew
rlabel metal1 s 11359 5623 11359 5623 4 dout_9
port 12 nsew
rlabel metal1 s 3871 5623 3871 5623 4 dout_3
port 6 nsew
rlabel metal1 s 6367 5623 6367 5623 4 dout_5
port 8 nsew
rlabel metal1 s 8863 5623 8863 5623 4 dout_7
port 10 nsew
rlabel metal1 s 12607 5623 12607 5623 4 dout_10
port 13 nsew
rlabel metal1 s 16351 5623 16351 5623 4 dout_13
port 16 nsew
rlabel metal1 s 20095 5623 20095 5623 4 dout_16
port 19 nsew
rlabel metal1 s 127 5623 127 5623 4 dout_0
port 3 nsew
rlabel metal1 s 2623 5623 2623 5623 4 dout_2
port 5 nsew
rlabel metal1 s 5119 5623 5119 5623 4 dout_4
port 7 nsew
rlabel metal1 s 18847 5623 18847 5623 4 dout_15
port 18 nsew
rlabel metal1 s 7615 5623 7615 5623 4 dout_6
port 9 nsew
rlabel metal1 s 17599 5623 17599 5623 4 dout_14
port 17 nsew
rlabel metal1 s 1375 5623 1375 5623 4 dout_1
port 4 nsew
rlabel metal1 s 13855 5623 13855 5623 4 dout_11
port 14 nsew
rlabel metal1 s 10111 5623 10111 5623 4 dout_8
port 11 nsew
rlabel metal1 s 14432 629 14432 629 4 br_23
port 218 nsew
rlabel metal1 s 12400 629 12400 629 4 bl_19
port 209 nsew
rlabel metal1 s 5072 629 5072 629 4 bl_8
port 187 nsew
rlabel metal1 s 6320 629 6320 629 4 bl_10
port 191 nsew
rlabel metal1 s 13808 629 13808 629 4 bl_22
port 215 nsew
rlabel metal1 s 11152 629 11152 629 4 bl_17
port 205 nsew
rlabel metal1 s 3824 629 3824 629 4 bl_6
port 183 nsew
rlabel metal1 s 704 629 704 629 4 br_1
port 174 nsew
rlabel metal1 s 19424 629 19424 629 4 br_31
port 234 nsew
rlabel metal1 s 13648 629 13648 629 4 bl_21
port 213 nsew
rlabel metal1 s 6784 629 6784 629 4 br_10
port 192 nsew
rlabel metal1 s 16768 629 16768 629 4 br_26
port 224 nsew
rlabel metal1 s 18016 629 18016 629 4 br_28
port 228 nsew
rlabel metal1 s 1168 629 1168 629 4 bl_1
port 173 nsew
rlabel metal1 s 16304 629 16304 629 4 bl_26
port 223 nsew
rlabel metal1 s 18640 629 18640 629 4 bl_29
port 229 nsew
rlabel metal1 s 15056 629 15056 629 4 bl_24
port 219 nsew
rlabel metal1 s 13024 629 13024 629 4 br_20
port 212 nsew
rlabel metal1 s 20048 629 20048 629 4 bl_32
port 235 nsew
rlabel metal1 s 19264 629 19264 629 4 br_30
port 232 nsew
rlabel metal1 s 14896 629 14896 629 4 bl_23
port 217 nsew
rlabel metal1 s 3040 629 3040 629 4 br_4
port 180 nsew
rlabel metal1 s 10688 629 10688 629 4 br_17
port 206 nsew
rlabel metal1 s 5536 629 5536 629 4 br_8
port 188 nsew
rlabel metal1 s 8816 629 8816 629 4 bl_14
port 199 nsew
rlabel metal1 s 12560 629 12560 629 4 bl_20
port 211 nsew
rlabel metal1 s 4912 629 4912 629 4 bl_7
port 185 nsew
rlabel metal1 s 10064 629 10064 629 4 bl_16
port 203 nsew
rlabel metal1 s 13184 629 13184 629 4 br_21
port 214 nsew
rlabel metal1 s 3664 629 3664 629 4 bl_5
port 181 nsew
rlabel metal1 s 4288 629 4288 629 4 br_6
port 184 nsew
rlabel metal1 s 16144 629 16144 629 4 bl_25
port 221 nsew
rlabel metal1 s 7408 629 7408 629 4 bl_11
port 193 nsew
rlabel metal1 s 6944 629 6944 629 4 br_11
port 194 nsew
rlabel metal1 s 9280 629 9280 629 4 br_14
port 200 nsew
rlabel metal1 s 8656 629 8656 629 4 bl_13
port 197 nsew
rlabel metal1 s 19888 629 19888 629 4 bl_31
port 233 nsew
rlabel metal1 s 15680 629 15680 629 4 br_25
port 222 nsew
rlabel metal1 s 9440 629 9440 629 4 br_15
port 202 nsew
rlabel metal1 s 3200 629 3200 629 4 br_5
port 182 nsew
rlabel metal1 s 11936 629 11936 629 4 br_19
port 210 nsew
rlabel metal1 s 9904 629 9904 629 4 bl_15
port 201 nsew
rlabel metal1 s 6160 629 6160 629 4 bl_9
port 189 nsew
rlabel metal1 s 17552 629 17552 629 4 bl_28
port 227 nsew
rlabel metal1 s 16928 629 16928 629 4 br_27
port 226 nsew
rlabel metal1 s 18800 629 18800 629 4 bl_30
port 231 nsew
rlabel metal1 s 1328 629 1328 629 4 bl_2
port 175 nsew
rlabel metal1 s 8032 629 8032 629 4 br_12
port 196 nsew
rlabel metal1 s 80 629 80 629 4 bl_0
port 171 nsew
rlabel metal1 s 2416 629 2416 629 4 bl_3
port 177 nsew
rlabel metal1 s 544 629 544 629 4 br_0
port 172 nsew
rlabel metal1 s 1792 629 1792 629 4 br_2
port 176 nsew
rlabel metal1 s 4448 629 4448 629 4 br_7
port 186 nsew
rlabel metal1 s 15520 629 15520 629 4 br_24
port 220 nsew
rlabel metal1 s 11312 629 11312 629 4 bl_18
port 207 nsew
rlabel metal1 s 18176 629 18176 629 4 br_29
port 230 nsew
rlabel metal1 s 7568 629 7568 629 4 bl_12
port 195 nsew
rlabel metal1 s 8192 629 8192 629 4 br_13
port 198 nsew
rlabel metal1 s 5696 629 5696 629 4 br_9
port 190 nsew
rlabel metal1 s 14272 629 14272 629 4 br_22
port 216 nsew
rlabel metal1 s 17392 629 17392 629 4 bl_27
port 225 nsew
rlabel metal1 s 11776 629 11776 629 4 br_18
port 208 nsew
rlabel metal1 s 2576 629 2576 629 4 bl_4
port 179 nsew
rlabel metal1 s 10528 629 10528 629 4 br_16
port 204 nsew
rlabel metal1 s 1952 629 1952 629 4 br_3
port 178 nsew
rlabel metal1 s 36112 629 36112 629 4 bl_57
port 285 nsew
rlabel metal1 s 36736 629 36736 629 4 br_58
port 288 nsew
rlabel metal1 s 29872 629 29872 629 4 bl_47
port 265 nsew
rlabel metal1 s 32368 629 32368 629 4 bl_51
port 273 nsew
rlabel metal1 s 30032 629 30032 629 4 bl_48
port 267 nsew
rlabel metal1 s 26912 629 26912 629 4 br_43
port 258 nsew
rlabel metal1 s 27376 629 27376 629 4 bl_43
port 257 nsew
rlabel metal1 s 24880 629 24880 629 4 bl_39
port 249 nsew
rlabel metal1 s 30656 629 30656 629 4 br_49
port 270 nsew
rlabel metal1 s 25504 629 25504 629 4 br_40
port 252 nsew
rlabel metal1 s 39856 629 39856 629 4 bl_63
port 297 nsew
rlabel metal1 s 39232 629 39232 629 4 br_62
port 296 nsew
rlabel metal1 s 34240 629 34240 629 4 br_54
port 280 nsew
rlabel metal1 s 25664 629 25664 629 4 br_41
port 254 nsew
rlabel metal1 s 28160 629 28160 629 4 br_45
port 262 nsew
rlabel metal1 s 27536 629 27536 629 4 bl_44
port 259 nsew
rlabel metal1 s 26752 629 26752 629 4 br_42
port 256 nsew
rlabel metal1 s 24256 629 24256 629 4 br_38
port 248 nsew
rlabel metal1 s 20512 629 20512 629 4 br_32
port 236 nsew
rlabel metal1 s 22544 629 22544 629 4 bl_36
port 243 nsew
rlabel metal1 s 26288 629 26288 629 4 bl_42
port 255 nsew
rlabel metal1 s 35488 629 35488 629 4 br_56
port 284 nsew
rlabel metal1 s 40480 629 40480 629 4 rbl_br
port 2 nsew
rlabel metal1 s 23632 629 23632 629 4 bl_37
port 245 nsew
rlabel metal1 s 39392 629 39392 629 4 br_63
port 298 nsew
rlabel metal1 s 23168 629 23168 629 4 br_37
port 246 nsew
rlabel metal1 s 30496 629 30496 629 4 br_48
port 268 nsew
rlabel metal1 s 29408 629 29408 629 4 br_47
port 266 nsew
rlabel metal1 s 23008 629 23008 629 4 br_36
port 244 nsew
rlabel metal1 s 32992 629 32992 629 4 br_52
port 276 nsew
rlabel metal1 s 28000 629 28000 629 4 br_44
port 260 nsew
rlabel metal1 s 28784 629 28784 629 4 bl_46
port 263 nsew
rlabel metal1 s 38768 629 38768 629 4 bl_62
port 295 nsew
rlabel metal1 s 25040 629 25040 629 4 bl_40
port 251 nsew
rlabel metal1 s 23792 629 23792 629 4 bl_38
port 247 nsew
rlabel metal1 s 21760 629 21760 629 4 br_34
port 240 nsew
rlabel metal1 s 37360 629 37360 629 4 bl_59
port 289 nsew
rlabel metal1 s 38608 629 38608 629 4 bl_61
port 293 nsew
rlabel metal1 s 40016 629 40016 629 4 rbl_bl
port 1 nsew
rlabel metal1 s 31904 629 31904 629 4 br_51
port 274 nsew
rlabel metal1 s 21296 629 21296 629 4 bl_34
port 239 nsew
rlabel metal1 s 24416 629 24416 629 4 br_39
port 250 nsew
rlabel metal1 s 32528 629 32528 629 4 bl_52
port 275 nsew
rlabel metal1 s 33616 629 33616 629 4 bl_53
port 277 nsew
rlabel metal1 s 26128 629 26128 629 4 bl_41
port 253 nsew
rlabel metal1 s 33152 629 33152 629 4 br_53
port 278 nsew
rlabel metal1 s 36896 629 36896 629 4 br_59
port 290 nsew
rlabel metal1 s 28624 629 28624 629 4 bl_45
port 261 nsew
rlabel metal1 s 20672 629 20672 629 4 br_33
port 238 nsew
rlabel metal1 s 38144 629 38144 629 4 br_61
port 294 nsew
rlabel metal1 s 21920 629 21920 629 4 br_35
port 242 nsew
rlabel metal1 s 36272 629 36272 629 4 bl_58
port 287 nsew
rlabel metal1 s 29248 629 29248 629 4 br_46
port 264 nsew
rlabel metal1 s 35648 629 35648 629 4 br_57
port 286 nsew
rlabel metal1 s 34400 629 34400 629 4 br_55
port 282 nsew
rlabel metal1 s 21136 629 21136 629 4 bl_33
port 237 nsew
rlabel metal1 s 34864 629 34864 629 4 bl_55
port 281 nsew
rlabel metal1 s 31744 629 31744 629 4 br_50
port 272 nsew
rlabel metal1 s 37984 629 37984 629 4 br_60
port 292 nsew
rlabel metal1 s 31280 629 31280 629 4 bl_50
port 271 nsew
rlabel metal1 s 31120 629 31120 629 4 bl_49
port 269 nsew
rlabel metal1 s 35024 629 35024 629 4 bl_56
port 283 nsew
rlabel metal1 s 22384 629 22384 629 4 bl_35
port 241 nsew
rlabel metal1 s 37520 629 37520 629 4 bl_60
port 291 nsew
rlabel metal1 s 33776 629 33776 629 4 bl_54
port 279 nsew
rlabel metal3 s 36573 5320 36573 5320 4 vdd
port 39 nsew
rlabel metal3 s 37809 4482 37809 4482 4 vdd
port 39 nsew
rlabel metal3 s 35325 5320 35325 5320 4 vdd
port 39 nsew
rlabel metal3 s 26589 5320 26589 5320 4 vdd
port 39 nsew
rlabel metal3 s 34065 4482 34065 4482 4 vdd
port 39 nsew
rlabel metal3 s 31581 5320 31581 5320 4 vdd
port 39 nsew
rlabel metal3 s 25341 5320 25341 5320 4 vdd
port 39 nsew
rlabel metal3 s 30333 5320 30333 5320 4 vdd
port 39 nsew
rlabel metal3 s 22833 4482 22833 4482 4 vdd
port 39 nsew
rlabel metal3 s 20349 5320 20349 5320 4 vdd
port 39 nsew
rlabel metal3 s 21585 4482 21585 4482 4 vdd
port 39 nsew
rlabel metal3 s 25329 4482 25329 4482 4 vdd
port 39 nsew
rlabel metal3 s 39069 5320 39069 5320 4 vdd
port 39 nsew
rlabel metal3 s 24093 5320 24093 5320 4 vdd
port 39 nsew
rlabel metal3 s 27837 5320 27837 5320 4 vdd
port 39 nsew
rlabel metal3 s 21597 5320 21597 5320 4 vdd
port 39 nsew
rlabel metal3 s 35313 4482 35313 4482 4 vdd
port 39 nsew
rlabel metal3 s 32817 4482 32817 4482 4 vdd
port 39 nsew
rlabel metal3 s 20337 4482 20337 4482 4 vdd
port 39 nsew
rlabel metal3 s 32829 5320 32829 5320 4 vdd
port 39 nsew
rlabel metal3 s 34077 5320 34077 5320 4 vdd
port 39 nsew
rlabel metal3 s 29085 5320 29085 5320 4 vdd
port 39 nsew
rlabel metal3 s 27825 4482 27825 4482 4 vdd
port 39 nsew
rlabel metal3 s 31569 4482 31569 4482 4 vdd
port 39 nsew
rlabel metal3 s 22845 5320 22845 5320 4 vdd
port 39 nsew
rlabel metal3 s 36561 4482 36561 4482 4 vdd
port 39 nsew
rlabel metal3 s 37821 5320 37821 5320 4 vdd
port 39 nsew
rlabel metal3 s 26577 4482 26577 4482 4 vdd
port 39 nsew
rlabel metal3 s 24081 4482 24081 4482 4 vdd
port 39 nsew
rlabel metal3 s 39057 4482 39057 4482 4 vdd
port 39 nsew
rlabel metal3 s 29073 4482 29073 4482 4 vdd
port 39 nsew
rlabel metal3 s 30321 4482 30321 4482 4 vdd
port 39 nsew
rlabel metal3 s 37821 5642 37821 5642 4 gnd
port 40 nsew
rlabel metal3 s 39139 3708 39139 3708 4 gnd
port 40 nsew
rlabel metal3 s 34147 3708 34147 3708 4 gnd
port 40 nsew
rlabel metal3 s 20349 5642 20349 5642 4 gnd
port 40 nsew
rlabel metal3 s 25341 5642 25341 5642 4 gnd
port 40 nsew
rlabel metal3 s 36643 3708 36643 3708 4 gnd
port 40 nsew
rlabel metal3 s 36573 5642 36573 5642 4 gnd
port 40 nsew
rlabel metal3 s 32899 3708 32899 3708 4 gnd
port 40 nsew
rlabel metal3 s 34077 5642 34077 5642 4 gnd
port 40 nsew
rlabel metal3 s 32829 5642 32829 5642 4 gnd
port 40 nsew
rlabel metal3 s 35325 5642 35325 5642 4 gnd
port 40 nsew
rlabel metal3 s 24163 3708 24163 3708 4 gnd
port 40 nsew
rlabel metal3 s 21667 3708 21667 3708 4 gnd
port 40 nsew
rlabel metal3 s 25411 3708 25411 3708 4 gnd
port 40 nsew
rlabel metal3 s 35395 3708 35395 3708 4 gnd
port 40 nsew
rlabel metal3 s 29155 3708 29155 3708 4 gnd
port 40 nsew
rlabel metal3 s 21597 5642 21597 5642 4 gnd
port 40 nsew
rlabel metal3 s 37891 3708 37891 3708 4 gnd
port 40 nsew
rlabel metal3 s 22845 5642 22845 5642 4 gnd
port 40 nsew
rlabel metal3 s 26659 3708 26659 3708 4 gnd
port 40 nsew
rlabel metal3 s 31651 3708 31651 3708 4 gnd
port 40 nsew
rlabel metal3 s 22915 3708 22915 3708 4 gnd
port 40 nsew
rlabel metal3 s 24093 5642 24093 5642 4 gnd
port 40 nsew
rlabel metal3 s 30333 5642 30333 5642 4 gnd
port 40 nsew
rlabel metal3 s 26589 5642 26589 5642 4 gnd
port 40 nsew
rlabel metal3 s 30403 3708 30403 3708 4 gnd
port 40 nsew
rlabel metal3 s 20419 3708 20419 3708 4 gnd
port 40 nsew
rlabel metal3 s 31581 5642 31581 5642 4 gnd
port 40 nsew
rlabel metal3 s 29085 5642 29085 5642 4 gnd
port 40 nsew
rlabel metal3 s 27837 5642 27837 5642 4 gnd
port 40 nsew
rlabel metal3 s 27907 3708 27907 3708 4 gnd
port 40 nsew
rlabel metal3 s 39069 5642 39069 5642 4 gnd
port 40 nsew
rlabel metal3 s 28080 1935 28080 1935 4 gnd
port 40 nsew
rlabel metal3 s 26832 1935 26832 1935 4 gnd
port 40 nsew
rlabel metal3 s 20592 1935 20592 1935 4 gnd
port 40 nsew
rlabel metal3 s 31824 1935 31824 1935 4 gnd
port 40 nsew
rlabel metal3 s 23088 1935 23088 1935 4 gnd
port 40 nsew
rlabel metal3 s 34320 1935 34320 1935 4 gnd
port 40 nsew
rlabel metal3 s 24336 1935 24336 1935 4 gnd
port 40 nsew
rlabel metal3 s 20280 981 20280 981 4 p_en_bar
port 38 nsew
rlabel metal3 s 38064 1935 38064 1935 4 gnd
port 40 nsew
rlabel metal3 s 25584 1935 25584 1935 4 gnd
port 40 nsew
rlabel metal3 s 39312 1935 39312 1935 4 gnd
port 40 nsew
rlabel metal3 s 35568 1935 35568 1935 4 gnd
port 40 nsew
rlabel metal3 s 21840 1935 21840 1935 4 gnd
port 40 nsew
rlabel metal3 s 36816 1935 36816 1935 4 gnd
port 40 nsew
rlabel metal3 s 33072 1935 33072 1935 4 gnd
port 40 nsew
rlabel metal3 s 30576 1935 30576 1935 4 gnd
port 40 nsew
rlabel metal3 s 29328 1935 29328 1935 4 gnd
port 40 nsew
rlabel metal3 s 4113 4482 4113 4482 4 vdd
port 39 nsew
rlabel metal3 s 16675 3708 16675 3708 4 gnd
port 40 nsew
rlabel metal3 s 4195 3708 4195 3708 4 gnd
port 40 nsew
rlabel metal3 s 16605 5642 16605 5642 4 gnd
port 40 nsew
rlabel metal3 s 2947 3708 2947 3708 4 gnd
port 40 nsew
rlabel metal3 s 7939 3708 7939 3708 4 gnd
port 40 nsew
rlabel metal3 s 5373 5642 5373 5642 4 gnd
port 40 nsew
rlabel metal3 s 19171 3708 19171 3708 4 gnd
port 40 nsew
rlabel metal3 s 10435 3708 10435 3708 4 gnd
port 40 nsew
rlabel metal3 s 19101 5320 19101 5320 4 vdd
port 39 nsew
rlabel metal3 s 19101 5642 19101 5642 4 gnd
port 40 nsew
rlabel metal3 s 10365 5320 10365 5320 4 vdd
port 39 nsew
rlabel metal3 s 4125 5320 4125 5320 4 vdd
port 39 nsew
rlabel metal3 s 17841 4482 17841 4482 4 vdd
port 39 nsew
rlabel metal3 s 381 5320 381 5320 4 vdd
port 39 nsew
rlabel metal3 s 17853 5642 17853 5642 4 gnd
port 40 nsew
rlabel metal3 s 9187 3708 9187 3708 4 gnd
port 40 nsew
rlabel metal3 s 14179 3708 14179 3708 4 gnd
port 40 nsew
rlabel metal3 s 15357 5642 15357 5642 4 gnd
port 40 nsew
rlabel metal3 s 16605 5320 16605 5320 4 vdd
port 39 nsew
rlabel metal3 s 12849 4482 12849 4482 4 vdd
port 39 nsew
rlabel metal3 s 17923 3708 17923 3708 4 gnd
port 40 nsew
rlabel metal3 s 2877 5320 2877 5320 4 vdd
port 39 nsew
rlabel metal3 s 9117 5320 9117 5320 4 vdd
port 39 nsew
rlabel metal3 s 11683 3708 11683 3708 4 gnd
port 40 nsew
rlabel metal3 s 15427 3708 15427 3708 4 gnd
port 40 nsew
rlabel metal3 s 5373 5320 5373 5320 4 vdd
port 39 nsew
rlabel metal3 s 12931 3708 12931 3708 4 gnd
port 40 nsew
rlabel metal3 s 12861 5320 12861 5320 4 vdd
port 39 nsew
rlabel metal3 s 6621 5642 6621 5642 4 gnd
port 40 nsew
rlabel metal3 s 7869 5320 7869 5320 4 vdd
port 39 nsew
rlabel metal3 s 2877 5642 2877 5642 4 gnd
port 40 nsew
rlabel metal3 s 381 5642 381 5642 4 gnd
port 40 nsew
rlabel metal3 s 451 3708 451 3708 4 gnd
port 40 nsew
rlabel metal3 s 11613 5642 11613 5642 4 gnd
port 40 nsew
rlabel metal3 s 11613 5320 11613 5320 4 vdd
port 39 nsew
rlabel metal3 s 7857 4482 7857 4482 4 vdd
port 39 nsew
rlabel metal3 s 16593 4482 16593 4482 4 vdd
port 39 nsew
rlabel metal3 s 14109 5320 14109 5320 4 vdd
port 39 nsew
rlabel metal3 s 4125 5642 4125 5642 4 gnd
port 40 nsew
rlabel metal3 s 14097 4482 14097 4482 4 vdd
port 39 nsew
rlabel metal3 s 10353 4482 10353 4482 4 vdd
port 39 nsew
rlabel metal3 s 19089 4482 19089 4482 4 vdd
port 39 nsew
rlabel metal3 s 6691 3708 6691 3708 4 gnd
port 40 nsew
rlabel metal3 s 15345 4482 15345 4482 4 vdd
port 39 nsew
rlabel metal3 s 19968 3556 19968 3556 4 s_en
port 37 nsew
rlabel metal3 s 5443 3708 5443 3708 4 gnd
port 40 nsew
rlabel metal3 s 12861 5642 12861 5642 4 gnd
port 40 nsew
rlabel metal3 s 19968 2840 19968 2840 4 sel_0
port 35 nsew
rlabel metal3 s 9360 1935 9360 1935 4 gnd
port 40 nsew
rlabel metal3 s 8112 1935 8112 1935 4 gnd
port 40 nsew
rlabel metal3 s 13104 1935 13104 1935 4 gnd
port 40 nsew
rlabel metal3 s 16848 1935 16848 1935 4 gnd
port 40 nsew
rlabel metal3 s 19344 1935 19344 1935 4 gnd
port 40 nsew
rlabel metal3 s 4368 1935 4368 1935 4 gnd
port 40 nsew
rlabel metal3 s 5616 1935 5616 1935 4 gnd
port 40 nsew
rlabel metal3 s 1872 1935 1872 1935 4 gnd
port 40 nsew
rlabel metal3 s 11856 1935 11856 1935 4 gnd
port 40 nsew
rlabel metal3 s 14352 1935 14352 1935 4 gnd
port 40 nsew
rlabel metal3 s 18096 1935 18096 1935 4 gnd
port 40 nsew
rlabel metal3 s 3120 1935 3120 1935 4 gnd
port 40 nsew
rlabel metal3 s 6864 1935 6864 1935 4 gnd
port 40 nsew
rlabel metal3 s 15600 1935 15600 1935 4 gnd
port 40 nsew
rlabel metal3 s 10608 1935 10608 1935 4 gnd
port 40 nsew
rlabel metal3 s 624 1935 624 1935 4 gnd
port 40 nsew
rlabel metal3 s 19968 2716 19968 2716 4 sel_1
port 36 nsew
rlabel metal3 s 6621 5320 6621 5320 4 vdd
port 39 nsew
rlabel metal3 s 14109 5642 14109 5642 4 gnd
port 40 nsew
rlabel metal3 s 369 4482 369 4482 4 vdd
port 39 nsew
rlabel metal3 s 6609 4482 6609 4482 4 vdd
port 39 nsew
rlabel metal3 s 10365 5642 10365 5642 4 gnd
port 40 nsew
rlabel metal3 s 1699 3708 1699 3708 4 gnd
port 40 nsew
rlabel metal3 s 1617 4482 1617 4482 4 vdd
port 39 nsew
rlabel metal3 s 17853 5320 17853 5320 4 vdd
port 39 nsew
rlabel metal3 s 9105 4482 9105 4482 4 vdd
port 39 nsew
rlabel metal3 s 1629 5320 1629 5320 4 vdd
port 39 nsew
rlabel metal3 s 7869 5642 7869 5642 4 gnd
port 40 nsew
rlabel metal3 s 11601 4482 11601 4482 4 vdd
port 39 nsew
rlabel metal3 s 9117 5642 9117 5642 4 gnd
port 40 nsew
rlabel metal3 s 2865 4482 2865 4482 4 vdd
port 39 nsew
rlabel metal3 s 15357 5320 15357 5320 4 vdd
port 39 nsew
rlabel metal3 s 5361 4482 5361 4482 4 vdd
port 39 nsew
rlabel metal3 s 1629 5642 1629 5642 4 gnd
port 40 nsew
rlabel metal3 s 5185 362 5185 362 4 vdd
port 39 nsew
rlabel metal3 s 1441 362 1441 362 4 vdd
port 39 nsew
rlabel metal3 s 8929 362 8929 362 4 vdd
port 39 nsew
rlabel metal3 s 15169 362 15169 362 4 vdd
port 39 nsew
rlabel metal3 s 13921 362 13921 362 4 vdd
port 39 nsew
rlabel metal3 s 16417 362 16417 362 4 vdd
port 39 nsew
rlabel metal3 s 17665 362 17665 362 4 vdd
port 39 nsew
rlabel metal3 s 17279 362 17279 362 4 vdd
port 39 nsew
rlabel metal3 s 18527 362 18527 362 4 vdd
port 39 nsew
rlabel metal3 s 13535 362 13535 362 4 vdd
port 39 nsew
rlabel metal3 s 14783 362 14783 362 4 vdd
port 39 nsew
rlabel metal3 s 2689 362 2689 362 4 vdd
port 39 nsew
rlabel metal3 s 19775 362 19775 362 4 vdd
port 39 nsew
rlabel metal3 s 2303 362 2303 362 4 vdd
port 39 nsew
rlabel metal3 s 18913 362 18913 362 4 vdd
port 39 nsew
rlabel metal3 s 8543 362 8543 362 4 vdd
port 39 nsew
rlabel metal3 s 11039 362 11039 362 4 vdd
port 39 nsew
rlabel metal3 s 4799 362 4799 362 4 vdd
port 39 nsew
rlabel metal3 s 12287 362 12287 362 4 vdd
port 39 nsew
rlabel metal3 s 7295 362 7295 362 4 vdd
port 39 nsew
rlabel metal3 s 3937 362 3937 362 4 vdd
port 39 nsew
rlabel metal3 s 6047 362 6047 362 4 vdd
port 39 nsew
rlabel metal3 s 10177 362 10177 362 4 vdd
port 39 nsew
rlabel metal3 s 1055 362 1055 362 4 vdd
port 39 nsew
rlabel metal3 s 193 362 193 362 4 vdd
port 39 nsew
rlabel metal3 s 9791 362 9791 362 4 vdd
port 39 nsew
rlabel metal3 s 7681 362 7681 362 4 vdd
port 39 nsew
rlabel metal3 s 3551 362 3551 362 4 vdd
port 39 nsew
rlabel metal3 s 16031 362 16031 362 4 vdd
port 39 nsew
rlabel metal3 s 20161 362 20161 362 4 vdd
port 39 nsew
rlabel metal3 s 11425 362 11425 362 4 vdd
port 39 nsew
rlabel metal3 s 6433 362 6433 362 4 vdd
port 39 nsew
rlabel metal3 s 12673 362 12673 362 4 vdd
port 39 nsew
rlabel metal3 s 32255 362 32255 362 4 vdd
port 39 nsew
rlabel metal3 s 27649 362 27649 362 4 vdd
port 39 nsew
rlabel metal3 s 21023 362 21023 362 4 vdd
port 39 nsew
rlabel metal3 s 27263 362 27263 362 4 vdd
port 39 nsew
rlabel metal3 s 37633 362 37633 362 4 vdd
port 39 nsew
rlabel metal3 s 24767 362 24767 362 4 vdd
port 39 nsew
rlabel metal3 s 36385 362 36385 362 4 vdd
port 39 nsew
rlabel metal3 s 21409 362 21409 362 4 vdd
port 39 nsew
rlabel metal3 s 34751 362 34751 362 4 vdd
port 39 nsew
rlabel metal3 s 31393 362 31393 362 4 vdd
port 39 nsew
rlabel metal3 s 35999 362 35999 362 4 vdd
port 39 nsew
rlabel metal3 s 38881 362 38881 362 4 vdd
port 39 nsew
rlabel metal3 s 23519 362 23519 362 4 vdd
port 39 nsew
rlabel metal3 s 39743 362 39743 362 4 vdd
port 39 nsew
rlabel metal3 s 25153 362 25153 362 4 vdd
port 39 nsew
rlabel metal3 s 32641 362 32641 362 4 vdd
port 39 nsew
rlabel metal3 s 26015 362 26015 362 4 vdd
port 39 nsew
rlabel metal3 s 40129 362 40129 362 4 vdd
port 39 nsew
rlabel metal3 s 22657 362 22657 362 4 vdd
port 39 nsew
rlabel metal3 s 33889 362 33889 362 4 vdd
port 39 nsew
rlabel metal3 s 22271 362 22271 362 4 vdd
port 39 nsew
rlabel metal3 s 28897 362 28897 362 4 vdd
port 39 nsew
rlabel metal3 s 38495 362 38495 362 4 vdd
port 39 nsew
rlabel metal3 s 33503 362 33503 362 4 vdd
port 39 nsew
rlabel metal3 s 30145 362 30145 362 4 vdd
port 39 nsew
rlabel metal3 s 37247 362 37247 362 4 vdd
port 39 nsew
rlabel metal3 s 29759 362 29759 362 4 vdd
port 39 nsew
rlabel metal3 s 35137 362 35137 362 4 vdd
port 39 nsew
rlabel metal3 s 26401 362 26401 362 4 vdd
port 39 nsew
rlabel metal3 s 28511 362 28511 362 4 vdd
port 39 nsew
rlabel metal3 s 31007 362 31007 362 4 vdd
port 39 nsew
rlabel metal3 s 23905 362 23905 362 4 vdd
port 39 nsew
<< properties >>
string FIXED_BBOX 0 0 40560 5750
string GDS_END 4847788
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 4738022
<< end >>
