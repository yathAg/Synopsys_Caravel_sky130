magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 5 21 1558 203
rect 29 -17 63 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 419 47 449 177
rect 503 47 533 177
rect 587 47 617 177
rect 671 47 701 177
rect 755 47 785 177
rect 922 47 952 177
rect 1006 47 1036 177
rect 1114 47 1144 177
rect 1198 47 1228 177
rect 1282 47 1312 177
rect 1366 47 1396 177
rect 1450 47 1480 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 419 297 449 497
rect 503 297 533 497
rect 587 297 617 497
rect 671 297 701 497
rect 862 297 892 497
rect 946 297 976 497
rect 1030 297 1060 497
rect 1114 297 1144 497
rect 1198 297 1228 497
rect 1282 297 1312 497
rect 1366 297 1396 497
rect 1450 297 1480 497
<< ndiff >>
rect 31 161 83 177
rect 31 127 39 161
rect 73 127 83 161
rect 31 93 83 127
rect 31 59 39 93
rect 73 59 83 93
rect 31 47 83 59
rect 113 93 167 177
rect 113 59 123 93
rect 157 59 167 93
rect 113 47 167 59
rect 197 157 251 177
rect 197 123 207 157
rect 241 123 251 157
rect 197 89 251 123
rect 197 55 207 89
rect 241 55 251 89
rect 197 47 251 55
rect 281 93 335 177
rect 281 59 291 93
rect 325 59 335 93
rect 281 47 335 59
rect 365 157 419 177
rect 365 123 375 157
rect 409 123 419 157
rect 365 89 419 123
rect 365 55 375 89
rect 409 55 419 89
rect 365 47 419 55
rect 449 93 503 177
rect 449 59 459 93
rect 493 59 503 93
rect 449 47 503 59
rect 533 157 587 177
rect 533 123 543 157
rect 577 123 587 157
rect 533 89 587 123
rect 533 55 543 89
rect 577 55 587 89
rect 533 47 587 55
rect 617 93 671 177
rect 617 59 627 93
rect 661 59 671 93
rect 617 47 671 59
rect 701 157 755 177
rect 701 123 711 157
rect 745 123 755 157
rect 701 89 755 123
rect 701 55 711 89
rect 745 55 755 89
rect 701 47 755 55
rect 785 89 922 177
rect 785 55 810 89
rect 844 55 878 89
rect 912 55 922 89
rect 785 47 922 55
rect 952 129 1006 177
rect 952 95 962 129
rect 996 95 1006 129
rect 952 47 1006 95
rect 1036 89 1114 177
rect 1036 55 1058 89
rect 1092 55 1114 89
rect 1036 47 1114 55
rect 1144 129 1198 177
rect 1144 95 1154 129
rect 1188 95 1198 129
rect 1144 47 1198 95
rect 1228 169 1282 177
rect 1228 135 1238 169
rect 1272 135 1282 169
rect 1228 47 1282 135
rect 1312 89 1366 177
rect 1312 55 1322 89
rect 1356 55 1366 89
rect 1312 47 1366 55
rect 1396 169 1450 177
rect 1396 135 1406 169
rect 1440 135 1450 169
rect 1396 47 1450 135
rect 1480 161 1532 177
rect 1480 127 1490 161
rect 1524 127 1532 161
rect 1480 93 1532 127
rect 1480 59 1490 93
rect 1524 59 1532 93
rect 1480 47 1532 59
<< pdiff >>
rect 27 489 83 497
rect 27 455 39 489
rect 73 455 83 489
rect 27 421 83 455
rect 27 387 39 421
rect 73 387 83 421
rect 27 353 83 387
rect 27 319 39 353
rect 73 319 83 353
rect 27 297 83 319
rect 113 485 167 497
rect 113 451 123 485
rect 157 451 167 485
rect 113 297 167 451
rect 197 489 251 497
rect 197 455 207 489
rect 241 455 251 489
rect 197 421 251 455
rect 197 387 207 421
rect 241 387 251 421
rect 197 353 251 387
rect 197 319 207 353
rect 241 319 251 353
rect 197 297 251 319
rect 281 485 335 497
rect 281 451 291 485
rect 325 451 335 485
rect 281 297 335 451
rect 365 489 419 497
rect 365 455 375 489
rect 409 455 419 489
rect 365 421 419 455
rect 365 387 375 421
rect 409 387 419 421
rect 365 353 419 387
rect 365 319 375 353
rect 409 319 419 353
rect 365 297 419 319
rect 449 369 503 497
rect 449 335 459 369
rect 493 335 503 369
rect 449 297 503 335
rect 533 489 587 497
rect 533 455 543 489
rect 577 455 587 489
rect 533 421 587 455
rect 533 387 543 421
rect 577 387 587 421
rect 533 297 587 387
rect 617 369 671 497
rect 617 335 627 369
rect 661 335 671 369
rect 617 297 671 335
rect 701 489 757 497
rect 701 455 711 489
rect 745 455 757 489
rect 701 427 757 455
rect 701 297 751 427
rect 811 349 862 497
rect 805 339 862 349
rect 805 305 818 339
rect 852 305 862 339
rect 805 297 862 305
rect 892 475 946 497
rect 892 441 902 475
rect 936 441 946 475
rect 892 407 946 441
rect 892 373 902 407
rect 936 373 946 407
rect 892 297 946 373
rect 976 339 1030 497
rect 976 305 986 339
rect 1020 305 1030 339
rect 976 297 1030 305
rect 1060 475 1114 497
rect 1060 441 1070 475
rect 1104 441 1114 475
rect 1060 407 1114 441
rect 1060 373 1070 407
rect 1104 373 1114 407
rect 1060 297 1114 373
rect 1144 475 1198 497
rect 1144 441 1154 475
rect 1188 441 1198 475
rect 1144 407 1198 441
rect 1144 373 1154 407
rect 1188 373 1198 407
rect 1144 339 1198 373
rect 1144 305 1154 339
rect 1188 305 1198 339
rect 1144 297 1198 305
rect 1228 489 1282 497
rect 1228 455 1238 489
rect 1272 455 1282 489
rect 1228 421 1282 455
rect 1228 387 1238 421
rect 1272 387 1282 421
rect 1228 297 1282 387
rect 1312 475 1366 497
rect 1312 441 1322 475
rect 1356 441 1366 475
rect 1312 407 1366 441
rect 1312 373 1322 407
rect 1356 373 1366 407
rect 1312 339 1366 373
rect 1312 305 1322 339
rect 1356 305 1366 339
rect 1312 297 1366 305
rect 1396 489 1450 497
rect 1396 455 1406 489
rect 1440 455 1450 489
rect 1396 421 1450 455
rect 1396 387 1406 421
rect 1440 387 1450 421
rect 1396 297 1450 387
rect 1480 423 1532 497
rect 1480 389 1490 423
rect 1524 389 1532 423
rect 1480 355 1532 389
rect 1480 321 1490 355
rect 1524 321 1532 355
rect 1480 297 1532 321
<< ndiffc >>
rect 39 127 73 161
rect 39 59 73 93
rect 123 59 157 93
rect 207 123 241 157
rect 207 55 241 89
rect 291 59 325 93
rect 375 123 409 157
rect 375 55 409 89
rect 459 59 493 93
rect 543 123 577 157
rect 543 55 577 89
rect 627 59 661 93
rect 711 123 745 157
rect 711 55 745 89
rect 810 55 844 89
rect 878 55 912 89
rect 962 95 996 129
rect 1058 55 1092 89
rect 1154 95 1188 129
rect 1238 135 1272 169
rect 1322 55 1356 89
rect 1406 135 1440 169
rect 1490 127 1524 161
rect 1490 59 1524 93
<< pdiffc >>
rect 39 455 73 489
rect 39 387 73 421
rect 39 319 73 353
rect 123 451 157 485
rect 207 455 241 489
rect 207 387 241 421
rect 207 319 241 353
rect 291 451 325 485
rect 375 455 409 489
rect 375 387 409 421
rect 375 319 409 353
rect 459 335 493 369
rect 543 455 577 489
rect 543 387 577 421
rect 627 335 661 369
rect 711 455 745 489
rect 818 305 852 339
rect 902 441 936 475
rect 902 373 936 407
rect 986 305 1020 339
rect 1070 441 1104 475
rect 1070 373 1104 407
rect 1154 441 1188 475
rect 1154 373 1188 407
rect 1154 305 1188 339
rect 1238 455 1272 489
rect 1238 387 1272 421
rect 1322 441 1356 475
rect 1322 373 1356 407
rect 1322 305 1356 339
rect 1406 455 1440 489
rect 1406 387 1440 421
rect 1490 389 1524 423
rect 1490 321 1524 355
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 419 497 449 523
rect 503 497 533 523
rect 587 497 617 523
rect 671 497 701 523
rect 862 497 892 523
rect 946 497 976 523
rect 1030 497 1060 523
rect 1114 497 1144 523
rect 1198 497 1228 523
rect 1282 497 1312 523
rect 1366 497 1396 523
rect 1450 497 1480 523
rect 83 259 113 297
rect 167 259 197 297
rect 251 259 281 297
rect 335 259 365 297
rect 83 249 365 259
rect 83 215 102 249
rect 136 215 170 249
rect 204 215 238 249
rect 272 215 306 249
rect 340 215 365 249
rect 83 205 365 215
rect 83 177 113 205
rect 167 177 197 205
rect 251 177 281 205
rect 335 177 365 205
rect 419 259 449 297
rect 503 259 533 297
rect 587 259 617 297
rect 671 259 701 297
rect 862 259 892 297
rect 946 259 976 297
rect 1030 259 1060 297
rect 1114 259 1144 297
rect 419 249 701 259
rect 419 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 701 249
rect 419 205 701 215
rect 419 177 449 205
rect 503 177 533 205
rect 587 177 617 205
rect 671 177 701 205
rect 755 249 1144 259
rect 755 215 771 249
rect 805 215 839 249
rect 873 215 907 249
rect 941 215 975 249
rect 1009 215 1043 249
rect 1077 215 1144 249
rect 755 205 1144 215
rect 755 177 785 205
rect 922 177 952 205
rect 1006 177 1036 205
rect 1114 177 1144 205
rect 1198 259 1228 297
rect 1282 259 1312 297
rect 1366 259 1396 297
rect 1450 259 1480 297
rect 1198 249 1495 259
rect 1198 215 1309 249
rect 1343 215 1377 249
rect 1411 215 1445 249
rect 1479 215 1495 249
rect 1198 205 1495 215
rect 1198 177 1228 205
rect 1282 177 1312 205
rect 1366 177 1396 205
rect 1450 177 1480 205
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 419 21 449 47
rect 503 21 533 47
rect 587 21 617 47
rect 671 21 701 47
rect 755 21 785 47
rect 922 21 952 47
rect 1006 21 1036 47
rect 1114 21 1144 47
rect 1198 21 1228 47
rect 1282 21 1312 47
rect 1366 21 1396 47
rect 1450 21 1480 47
<< polycont >>
rect 102 215 136 249
rect 170 215 204 249
rect 238 215 272 249
rect 306 215 340 249
rect 435 215 469 249
rect 503 215 537 249
rect 571 215 605 249
rect 639 215 673 249
rect 771 215 805 249
rect 839 215 873 249
rect 907 215 941 249
rect 975 215 1009 249
rect 1043 215 1077 249
rect 1309 215 1343 249
rect 1377 215 1411 249
rect 1445 215 1479 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 489 89 493
rect 18 455 39 489
rect 73 455 89 489
rect 18 421 89 455
rect 18 387 39 421
rect 73 387 89 421
rect 123 485 157 527
rect 123 413 157 451
rect 191 489 257 493
rect 191 455 207 489
rect 241 455 257 489
rect 191 421 257 455
rect 18 379 89 387
rect 191 387 207 421
rect 241 387 257 421
rect 291 485 325 527
rect 291 413 325 451
rect 359 489 777 493
rect 359 455 375 489
rect 409 455 543 489
rect 577 455 711 489
rect 745 455 777 489
rect 359 441 777 455
rect 816 475 1120 493
rect 816 441 902 475
rect 936 441 1070 475
rect 1104 441 1120 475
rect 359 421 425 441
rect 191 379 257 387
rect 359 387 375 421
rect 409 387 425 421
rect 527 421 593 441
rect 359 379 425 387
rect 18 353 425 379
rect 18 319 39 353
rect 73 319 207 353
rect 241 319 375 353
rect 409 319 425 353
rect 459 369 493 407
rect 527 387 543 421
rect 577 387 593 421
rect 816 407 1120 441
rect 627 373 902 407
rect 936 373 1070 407
rect 1104 373 1120 407
rect 1154 475 1188 493
rect 1154 407 1188 441
rect 1222 489 1288 527
rect 1222 455 1238 489
rect 1272 455 1288 489
rect 1222 421 1288 455
rect 1222 387 1238 421
rect 1272 387 1288 421
rect 1222 378 1288 387
rect 1322 475 1356 493
rect 1322 407 1356 441
rect 627 369 721 373
rect 493 335 627 353
rect 661 335 721 369
rect 1154 339 1188 373
rect 1390 489 1456 527
rect 1390 455 1406 489
rect 1440 455 1456 489
rect 1390 421 1456 455
rect 1390 387 1406 421
rect 1440 387 1456 421
rect 1390 378 1456 387
rect 1490 423 1547 493
rect 1524 389 1547 423
rect 1322 339 1356 373
rect 1490 355 1547 389
rect 459 319 721 335
rect 755 305 818 339
rect 852 305 986 339
rect 1020 305 1154 339
rect 1188 305 1322 339
rect 1356 321 1490 339
rect 1524 321 1547 355
rect 1356 305 1547 321
rect 755 289 1547 305
rect 18 249 356 285
rect 18 215 102 249
rect 136 215 170 249
rect 204 215 238 249
rect 272 215 306 249
rect 340 215 356 249
rect 18 211 356 215
rect 390 249 721 285
rect 390 215 435 249
rect 469 215 503 249
rect 537 215 571 249
rect 605 215 639 249
rect 673 215 721 249
rect 390 211 721 215
rect 755 249 1188 255
rect 755 215 771 249
rect 805 215 839 249
rect 873 215 907 249
rect 941 215 975 249
rect 1009 215 1043 249
rect 1077 215 1188 249
rect 755 211 1188 215
rect 1222 177 1259 289
rect 1293 249 1547 255
rect 1293 215 1309 249
rect 1343 215 1377 249
rect 1411 215 1445 249
rect 1479 215 1547 249
rect 1293 211 1547 215
rect 18 161 1188 177
rect 18 127 39 161
rect 73 157 1188 161
rect 73 143 207 157
rect 73 127 89 143
rect 18 93 89 127
rect 191 123 207 143
rect 241 143 375 157
rect 241 123 257 143
rect 18 59 39 93
rect 73 59 89 93
rect 18 51 89 59
rect 123 93 157 109
rect 123 17 157 59
rect 191 89 257 123
rect 359 123 375 143
rect 409 143 543 157
rect 409 123 425 143
rect 191 55 207 89
rect 241 55 257 89
rect 191 51 257 55
rect 291 93 325 109
rect 291 17 325 59
rect 359 89 425 123
rect 527 123 543 143
rect 577 143 711 157
rect 577 123 593 143
rect 359 55 375 89
rect 409 55 425 89
rect 359 51 425 55
rect 459 93 493 109
rect 459 17 493 59
rect 527 89 593 123
rect 695 123 711 143
rect 745 143 1188 157
rect 745 123 761 143
rect 527 55 543 89
rect 577 55 593 89
rect 527 51 593 55
rect 627 93 661 109
rect 627 17 661 59
rect 695 89 761 123
rect 962 129 996 143
rect 695 55 711 89
rect 745 55 761 89
rect 695 51 761 55
rect 799 89 928 109
rect 799 55 810 89
rect 844 55 878 89
rect 912 55 928 89
rect 1154 129 1188 143
rect 1222 169 1456 177
rect 1222 135 1238 169
rect 1272 135 1406 169
rect 1440 135 1456 169
rect 1222 129 1456 135
rect 1490 161 1547 177
rect 962 79 996 95
rect 1030 89 1120 109
rect 799 17 928 55
rect 1030 55 1058 89
rect 1092 55 1120 89
rect 1030 17 1120 55
rect 1524 127 1547 161
rect 1490 95 1547 127
rect 1154 93 1547 95
rect 1154 89 1490 93
rect 1154 55 1322 89
rect 1356 59 1490 89
rect 1524 59 1547 93
rect 1356 55 1547 59
rect 1154 51 1547 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 766 221 800 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 674 221 708 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 766 289 800 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 857 289 891 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 949 289 983 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1041 289 1075 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1133 289 1167 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1225 289 1259 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1317 289 1351 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1409 289 1443 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1501 289 1535 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1501 425 1535 459 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1501 357 1535 391 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1501 221 1535 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1409 221 1443 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1317 221 1351 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1225 153 1259 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1225 221 1259 255 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o31ai_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 1453680
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1439196
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 7.820 0.000 
<< end >>
