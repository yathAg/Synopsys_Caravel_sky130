magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< dnwell >>
rect -38 -38 1072 4993
<< nwell >>
rect -101 5076 121 12303
rect -118 4908 1119 5076
rect -118 168 168 4908
rect 782 168 1119 4908
rect -118 150 1119 168
rect -118 -134 1152 150
<< pwell >>
rect 228 228 722 4848
<< mvnmos >>
rect 415 3714 535 4714
rect 415 2593 535 3593
rect 415 1472 535 2472
rect 415 362 535 1362
<< mvndiff >>
rect 362 4702 415 4714
rect 362 4668 370 4702
rect 404 4668 415 4702
rect 362 4634 415 4668
rect 362 4600 370 4634
rect 404 4600 415 4634
rect 362 4566 415 4600
rect 362 4532 370 4566
rect 404 4532 415 4566
rect 362 4498 415 4532
rect 362 4464 370 4498
rect 404 4464 415 4498
rect 362 4430 415 4464
rect 362 4396 370 4430
rect 404 4396 415 4430
rect 362 4362 415 4396
rect 362 4328 370 4362
rect 404 4328 415 4362
rect 362 4294 415 4328
rect 362 4260 370 4294
rect 404 4260 415 4294
rect 362 4226 415 4260
rect 362 4192 370 4226
rect 404 4192 415 4226
rect 362 4158 415 4192
rect 362 4124 370 4158
rect 404 4124 415 4158
rect 362 4090 415 4124
rect 362 4056 370 4090
rect 404 4056 415 4090
rect 362 4022 415 4056
rect 362 3988 370 4022
rect 404 3988 415 4022
rect 362 3954 415 3988
rect 362 3920 370 3954
rect 404 3920 415 3954
rect 362 3886 415 3920
rect 362 3852 370 3886
rect 404 3852 415 3886
rect 362 3818 415 3852
rect 362 3784 370 3818
rect 404 3784 415 3818
rect 362 3714 415 3784
rect 535 4702 588 4714
rect 535 4668 546 4702
rect 580 4668 588 4702
rect 535 4634 588 4668
rect 535 4600 546 4634
rect 580 4600 588 4634
rect 535 4566 588 4600
rect 535 4532 546 4566
rect 580 4532 588 4566
rect 535 4498 588 4532
rect 535 4464 546 4498
rect 580 4464 588 4498
rect 535 4430 588 4464
rect 535 4396 546 4430
rect 580 4396 588 4430
rect 535 4362 588 4396
rect 535 4328 546 4362
rect 580 4328 588 4362
rect 535 4294 588 4328
rect 535 4260 546 4294
rect 580 4260 588 4294
rect 535 4226 588 4260
rect 535 4192 546 4226
rect 580 4192 588 4226
rect 535 4158 588 4192
rect 535 4124 546 4158
rect 580 4124 588 4158
rect 535 4090 588 4124
rect 535 4056 546 4090
rect 580 4056 588 4090
rect 535 4022 588 4056
rect 535 3988 546 4022
rect 580 3988 588 4022
rect 535 3954 588 3988
rect 535 3920 546 3954
rect 580 3920 588 3954
rect 535 3886 588 3920
rect 535 3852 546 3886
rect 580 3852 588 3886
rect 535 3818 588 3852
rect 535 3784 546 3818
rect 580 3784 588 3818
rect 535 3714 588 3784
rect 362 3581 415 3593
rect 362 3547 370 3581
rect 404 3547 415 3581
rect 362 3513 415 3547
rect 362 3479 370 3513
rect 404 3479 415 3513
rect 362 3445 415 3479
rect 362 3411 370 3445
rect 404 3411 415 3445
rect 362 3377 415 3411
rect 362 3343 370 3377
rect 404 3343 415 3377
rect 362 3309 415 3343
rect 362 3275 370 3309
rect 404 3275 415 3309
rect 362 3241 415 3275
rect 362 3207 370 3241
rect 404 3207 415 3241
rect 362 3173 415 3207
rect 362 3139 370 3173
rect 404 3139 415 3173
rect 362 3105 415 3139
rect 362 3071 370 3105
rect 404 3071 415 3105
rect 362 3037 415 3071
rect 362 3003 370 3037
rect 404 3003 415 3037
rect 362 2969 415 3003
rect 362 2935 370 2969
rect 404 2935 415 2969
rect 362 2901 415 2935
rect 362 2867 370 2901
rect 404 2867 415 2901
rect 362 2833 415 2867
rect 362 2799 370 2833
rect 404 2799 415 2833
rect 362 2765 415 2799
rect 362 2731 370 2765
rect 404 2731 415 2765
rect 362 2697 415 2731
rect 362 2663 370 2697
rect 404 2663 415 2697
rect 362 2593 415 2663
rect 535 3581 588 3593
rect 535 3547 546 3581
rect 580 3547 588 3581
rect 535 3513 588 3547
rect 535 3479 546 3513
rect 580 3479 588 3513
rect 535 3445 588 3479
rect 535 3411 546 3445
rect 580 3411 588 3445
rect 535 3377 588 3411
rect 535 3343 546 3377
rect 580 3343 588 3377
rect 535 3309 588 3343
rect 535 3275 546 3309
rect 580 3275 588 3309
rect 535 3241 588 3275
rect 535 3207 546 3241
rect 580 3207 588 3241
rect 535 3173 588 3207
rect 535 3139 546 3173
rect 580 3139 588 3173
rect 535 3105 588 3139
rect 535 3071 546 3105
rect 580 3071 588 3105
rect 535 3037 588 3071
rect 535 3003 546 3037
rect 580 3003 588 3037
rect 535 2969 588 3003
rect 535 2935 546 2969
rect 580 2935 588 2969
rect 535 2901 588 2935
rect 535 2867 546 2901
rect 580 2867 588 2901
rect 535 2833 588 2867
rect 535 2799 546 2833
rect 580 2799 588 2833
rect 535 2765 588 2799
rect 535 2731 546 2765
rect 580 2731 588 2765
rect 535 2697 588 2731
rect 535 2663 546 2697
rect 580 2663 588 2697
rect 535 2593 588 2663
rect 362 2460 415 2472
rect 362 2426 370 2460
rect 404 2426 415 2460
rect 362 2392 415 2426
rect 362 2358 370 2392
rect 404 2358 415 2392
rect 362 2324 415 2358
rect 362 2290 370 2324
rect 404 2290 415 2324
rect 362 2256 415 2290
rect 362 2222 370 2256
rect 404 2222 415 2256
rect 362 2188 415 2222
rect 362 2154 370 2188
rect 404 2154 415 2188
rect 362 2120 415 2154
rect 362 2086 370 2120
rect 404 2086 415 2120
rect 362 2052 415 2086
rect 362 2018 370 2052
rect 404 2018 415 2052
rect 362 1984 415 2018
rect 362 1950 370 1984
rect 404 1950 415 1984
rect 362 1916 415 1950
rect 362 1882 370 1916
rect 404 1882 415 1916
rect 362 1848 415 1882
rect 362 1814 370 1848
rect 404 1814 415 1848
rect 362 1780 415 1814
rect 362 1746 370 1780
rect 404 1746 415 1780
rect 362 1712 415 1746
rect 362 1678 370 1712
rect 404 1678 415 1712
rect 362 1644 415 1678
rect 362 1610 370 1644
rect 404 1610 415 1644
rect 362 1576 415 1610
rect 362 1542 370 1576
rect 404 1542 415 1576
rect 362 1472 415 1542
rect 535 2460 588 2472
rect 535 2426 546 2460
rect 580 2426 588 2460
rect 535 2392 588 2426
rect 535 2358 546 2392
rect 580 2358 588 2392
rect 535 2324 588 2358
rect 535 2290 546 2324
rect 580 2290 588 2324
rect 535 2256 588 2290
rect 535 2222 546 2256
rect 580 2222 588 2256
rect 535 2188 588 2222
rect 535 2154 546 2188
rect 580 2154 588 2188
rect 535 2120 588 2154
rect 535 2086 546 2120
rect 580 2086 588 2120
rect 535 2052 588 2086
rect 535 2018 546 2052
rect 580 2018 588 2052
rect 535 1984 588 2018
rect 535 1950 546 1984
rect 580 1950 588 1984
rect 535 1916 588 1950
rect 535 1882 546 1916
rect 580 1882 588 1916
rect 535 1848 588 1882
rect 535 1814 546 1848
rect 580 1814 588 1848
rect 535 1780 588 1814
rect 535 1746 546 1780
rect 580 1746 588 1780
rect 535 1712 588 1746
rect 535 1678 546 1712
rect 580 1678 588 1712
rect 535 1644 588 1678
rect 535 1610 546 1644
rect 580 1610 588 1644
rect 535 1576 588 1610
rect 535 1542 546 1576
rect 580 1542 588 1576
rect 535 1472 588 1542
rect 362 1292 415 1362
rect 362 1258 370 1292
rect 404 1258 415 1292
rect 362 1224 415 1258
rect 362 1190 370 1224
rect 404 1190 415 1224
rect 362 1156 415 1190
rect 362 1122 370 1156
rect 404 1122 415 1156
rect 362 1088 415 1122
rect 362 1054 370 1088
rect 404 1054 415 1088
rect 362 1020 415 1054
rect 362 986 370 1020
rect 404 986 415 1020
rect 362 952 415 986
rect 362 918 370 952
rect 404 918 415 952
rect 362 884 415 918
rect 362 850 370 884
rect 404 850 415 884
rect 362 816 415 850
rect 362 782 370 816
rect 404 782 415 816
rect 362 748 415 782
rect 362 714 370 748
rect 404 714 415 748
rect 362 680 415 714
rect 362 646 370 680
rect 404 646 415 680
rect 362 612 415 646
rect 362 578 370 612
rect 404 578 415 612
rect 362 544 415 578
rect 362 510 370 544
rect 404 510 415 544
rect 362 476 415 510
rect 362 442 370 476
rect 404 442 415 476
rect 362 408 415 442
rect 362 374 370 408
rect 404 374 415 408
rect 362 362 415 374
rect 535 1292 588 1362
rect 535 1258 546 1292
rect 580 1258 588 1292
rect 535 1224 588 1258
rect 535 1190 546 1224
rect 580 1190 588 1224
rect 535 1156 588 1190
rect 535 1122 546 1156
rect 580 1122 588 1156
rect 535 1088 588 1122
rect 535 1054 546 1088
rect 580 1054 588 1088
rect 535 1020 588 1054
rect 535 986 546 1020
rect 580 986 588 1020
rect 535 952 588 986
rect 535 918 546 952
rect 580 918 588 952
rect 535 884 588 918
rect 535 850 546 884
rect 580 850 588 884
rect 535 816 588 850
rect 535 782 546 816
rect 580 782 588 816
rect 535 748 588 782
rect 535 714 546 748
rect 580 714 588 748
rect 535 680 588 714
rect 535 646 546 680
rect 580 646 588 680
rect 535 612 588 646
rect 535 578 546 612
rect 580 578 588 612
rect 535 544 588 578
rect 535 510 546 544
rect 580 510 588 544
rect 535 476 588 510
rect 535 442 546 476
rect 580 442 588 476
rect 535 408 588 442
rect 535 374 546 408
rect 580 374 588 408
rect 535 362 588 374
<< mvndiffc >>
rect 370 4668 404 4702
rect 370 4600 404 4634
rect 370 4532 404 4566
rect 370 4464 404 4498
rect 370 4396 404 4430
rect 370 4328 404 4362
rect 370 4260 404 4294
rect 370 4192 404 4226
rect 370 4124 404 4158
rect 370 4056 404 4090
rect 370 3988 404 4022
rect 370 3920 404 3954
rect 370 3852 404 3886
rect 370 3784 404 3818
rect 546 4668 580 4702
rect 546 4600 580 4634
rect 546 4532 580 4566
rect 546 4464 580 4498
rect 546 4396 580 4430
rect 546 4328 580 4362
rect 546 4260 580 4294
rect 546 4192 580 4226
rect 546 4124 580 4158
rect 546 4056 580 4090
rect 546 3988 580 4022
rect 546 3920 580 3954
rect 546 3852 580 3886
rect 546 3784 580 3818
rect 370 3547 404 3581
rect 370 3479 404 3513
rect 370 3411 404 3445
rect 370 3343 404 3377
rect 370 3275 404 3309
rect 370 3207 404 3241
rect 370 3139 404 3173
rect 370 3071 404 3105
rect 370 3003 404 3037
rect 370 2935 404 2969
rect 370 2867 404 2901
rect 370 2799 404 2833
rect 370 2731 404 2765
rect 370 2663 404 2697
rect 546 3547 580 3581
rect 546 3479 580 3513
rect 546 3411 580 3445
rect 546 3343 580 3377
rect 546 3275 580 3309
rect 546 3207 580 3241
rect 546 3139 580 3173
rect 546 3071 580 3105
rect 546 3003 580 3037
rect 546 2935 580 2969
rect 546 2867 580 2901
rect 546 2799 580 2833
rect 546 2731 580 2765
rect 546 2663 580 2697
rect 370 2426 404 2460
rect 370 2358 404 2392
rect 370 2290 404 2324
rect 370 2222 404 2256
rect 370 2154 404 2188
rect 370 2086 404 2120
rect 370 2018 404 2052
rect 370 1950 404 1984
rect 370 1882 404 1916
rect 370 1814 404 1848
rect 370 1746 404 1780
rect 370 1678 404 1712
rect 370 1610 404 1644
rect 370 1542 404 1576
rect 546 2426 580 2460
rect 546 2358 580 2392
rect 546 2290 580 2324
rect 546 2222 580 2256
rect 546 2154 580 2188
rect 546 2086 580 2120
rect 546 2018 580 2052
rect 546 1950 580 1984
rect 546 1882 580 1916
rect 546 1814 580 1848
rect 546 1746 580 1780
rect 546 1678 580 1712
rect 546 1610 580 1644
rect 546 1542 580 1576
rect 370 1258 404 1292
rect 370 1190 404 1224
rect 370 1122 404 1156
rect 370 1054 404 1088
rect 370 986 404 1020
rect 370 918 404 952
rect 370 850 404 884
rect 370 782 404 816
rect 370 714 404 748
rect 370 646 404 680
rect 370 578 404 612
rect 370 510 404 544
rect 370 442 404 476
rect 370 374 404 408
rect 546 1258 580 1292
rect 546 1190 580 1224
rect 546 1122 580 1156
rect 546 1054 580 1088
rect 546 986 580 1020
rect 546 918 580 952
rect 546 850 580 884
rect 546 782 580 816
rect 546 714 580 748
rect 546 646 580 680
rect 546 578 580 612
rect 546 510 580 544
rect 546 442 580 476
rect 546 374 580 408
<< mvpsubdiff >>
rect 254 4788 278 4822
rect 312 4788 391 4822
rect 425 4788 525 4822
rect 559 4798 696 4822
rect 559 4788 662 4798
rect 254 4728 288 4788
rect 662 4729 696 4764
rect 254 4659 288 4694
rect 254 4590 288 4625
rect 254 4521 288 4556
rect 254 4452 288 4487
rect 254 4383 288 4418
rect 254 4314 288 4349
rect 254 4245 288 4280
rect 254 4176 288 4211
rect 254 4107 288 4142
rect 254 4038 288 4073
rect 254 3969 288 4004
rect 254 3900 288 3935
rect 254 3831 288 3866
rect 254 3762 288 3797
rect 254 3693 288 3728
rect 662 4660 696 4695
rect 662 4591 696 4626
rect 662 4522 696 4557
rect 662 4453 696 4488
rect 662 4384 696 4419
rect 662 4315 696 4350
rect 662 4246 696 4281
rect 662 4177 696 4212
rect 662 4108 696 4143
rect 662 4039 696 4074
rect 662 3970 696 4005
rect 662 3901 696 3936
rect 662 3832 696 3867
rect 662 3763 696 3798
rect 254 3624 288 3659
rect 662 3694 696 3729
rect 662 3625 696 3660
rect 254 3555 288 3590
rect 254 3486 288 3521
rect 254 3417 288 3452
rect 254 3348 288 3383
rect 254 3279 288 3314
rect 254 3210 288 3245
rect 254 3141 288 3176
rect 254 3072 288 3107
rect 254 3003 288 3038
rect 254 2934 288 2969
rect 254 2865 288 2900
rect 254 2796 288 2831
rect 254 2727 288 2762
rect 254 2658 288 2693
rect 254 2589 288 2624
rect 662 3556 696 3591
rect 662 3487 696 3522
rect 662 3418 696 3453
rect 662 3349 696 3384
rect 662 3280 696 3315
rect 662 3211 696 3246
rect 662 3142 696 3177
rect 662 3073 696 3108
rect 662 3004 696 3039
rect 662 2935 696 2970
rect 662 2866 696 2901
rect 662 2797 696 2832
rect 662 2728 696 2763
rect 662 2659 696 2694
rect 254 2520 288 2555
rect 254 2451 288 2486
rect 662 2590 696 2625
rect 662 2521 696 2556
rect 254 2382 288 2417
rect 254 2313 288 2348
rect 254 2244 288 2279
rect 254 2175 288 2210
rect 254 2106 288 2141
rect 254 2037 288 2072
rect 254 1968 288 2003
rect 254 1899 288 1934
rect 254 1830 288 1865
rect 254 1761 288 1796
rect 254 1692 288 1727
rect 254 1623 288 1658
rect 254 1554 288 1589
rect 254 1485 288 1520
rect 662 2452 696 2487
rect 662 2383 696 2418
rect 662 2314 696 2349
rect 662 2245 696 2280
rect 662 2176 696 2211
rect 662 2107 696 2142
rect 662 2038 696 2073
rect 662 1969 696 2004
rect 662 1900 696 1935
rect 662 1831 696 1866
rect 662 1762 696 1797
rect 662 1693 696 1728
rect 662 1624 696 1659
rect 662 1555 696 1590
rect 662 1486 696 1521
rect 254 1416 288 1451
rect 254 1347 288 1382
rect 662 1417 696 1452
rect 254 1278 288 1313
rect 254 1209 288 1244
rect 254 1140 288 1175
rect 254 1071 288 1106
rect 254 1002 288 1037
rect 254 933 288 968
rect 254 864 288 899
rect 254 795 288 830
rect 254 726 288 761
rect 254 657 288 692
rect 254 588 288 623
rect 254 519 288 554
rect 254 450 288 485
rect 254 381 288 416
rect 662 1348 696 1383
rect 662 1279 696 1314
rect 662 1210 696 1245
rect 662 1141 696 1176
rect 662 1072 696 1107
rect 662 1003 696 1038
rect 662 934 696 969
rect 662 865 696 900
rect 662 796 696 831
rect 662 727 696 762
rect 662 658 696 693
rect 662 589 696 624
rect 662 520 696 555
rect 662 451 696 486
rect 662 382 696 417
rect 254 312 288 347
rect 662 288 696 348
rect 288 278 352 288
rect 254 254 352 278
rect 386 254 423 288
rect 457 254 494 288
rect 528 254 566 288
rect 600 254 638 288
rect 672 254 696 288
<< mvnsubdiff >>
rect -35 12213 68 12237
rect -35 12179 -7 12213
rect 27 12179 68 12213
rect -35 12145 68 12179
rect -35 12111 -7 12145
rect 27 12111 68 12145
rect -35 12077 68 12111
rect -35 12043 -7 12077
rect 27 12043 68 12077
rect -35 12009 68 12043
rect -35 11975 -7 12009
rect 27 11975 68 12009
rect -35 11941 68 11975
rect -35 11907 -7 11941
rect 27 11907 68 11941
rect -35 11873 68 11907
rect -35 11839 -7 11873
rect 27 11839 68 11873
rect -35 11805 68 11839
rect -35 11771 -7 11805
rect 27 11771 68 11805
rect -35 11737 68 11771
rect -35 11703 -7 11737
rect 27 11703 68 11737
rect -35 11669 68 11703
rect -35 11635 -7 11669
rect 27 11635 68 11669
rect -35 11601 68 11635
rect -35 11567 -7 11601
rect 27 11567 68 11601
rect -35 11533 68 11567
rect -35 11499 -7 11533
rect 27 11499 68 11533
rect -35 11465 68 11499
rect -35 11431 -7 11465
rect 27 11431 68 11465
rect -35 11397 68 11431
rect -35 11363 -7 11397
rect 27 11363 68 11397
rect -35 11329 68 11363
rect -35 11295 -7 11329
rect 27 11295 68 11329
rect -35 11261 68 11295
rect -35 11227 -7 11261
rect 27 11227 68 11261
rect -35 11193 68 11227
rect -35 11159 -7 11193
rect 27 11159 68 11193
rect -35 11125 68 11159
rect -35 11091 -7 11125
rect 27 11091 68 11125
rect -35 11057 68 11091
rect -35 11023 -7 11057
rect 27 11023 68 11057
rect -35 10989 68 11023
rect -35 10955 -7 10989
rect 27 10955 68 10989
rect -35 10921 68 10955
rect -35 10887 -7 10921
rect 27 10887 68 10921
rect -35 10853 68 10887
rect -35 10819 -7 10853
rect 27 10819 68 10853
rect -35 10785 68 10819
rect -35 10751 -7 10785
rect 27 10751 68 10785
rect -35 10717 68 10751
rect -35 10683 -7 10717
rect 27 10683 68 10717
rect -35 10649 68 10683
rect -35 10615 -7 10649
rect 27 10615 68 10649
rect -35 10581 68 10615
rect -35 10547 -7 10581
rect 27 10547 68 10581
rect -35 10513 68 10547
rect -35 10479 -7 10513
rect 27 10479 68 10513
rect -35 10445 68 10479
rect -35 10411 -7 10445
rect 27 10411 68 10445
rect -35 10377 68 10411
rect -35 10343 -7 10377
rect 27 10343 68 10377
rect -35 10309 68 10343
rect -35 10275 -7 10309
rect 27 10275 68 10309
rect -35 10241 68 10275
rect -35 10207 -7 10241
rect 27 10207 68 10241
rect -35 10173 68 10207
rect -35 10139 -7 10173
rect 27 10139 68 10173
rect -35 10105 68 10139
rect -35 10071 -7 10105
rect 27 10071 68 10105
rect -35 10037 68 10071
rect -35 10003 -7 10037
rect 27 10003 68 10037
rect -35 9969 68 10003
rect -35 9935 -7 9969
rect 27 9935 68 9969
rect -35 9901 68 9935
rect -35 9867 -7 9901
rect 27 9867 68 9901
rect -35 9833 68 9867
rect -35 9799 -7 9833
rect 27 9799 68 9833
rect -35 9765 68 9799
rect -35 9731 -7 9765
rect 27 9731 68 9765
rect -35 9697 68 9731
rect -35 9663 -7 9697
rect 27 9663 68 9697
rect -35 9629 68 9663
rect -35 9595 -7 9629
rect 27 9595 68 9629
rect -35 9561 68 9595
rect -35 9527 -7 9561
rect 27 9527 68 9561
rect -35 9493 68 9527
rect -35 9459 -7 9493
rect 27 9459 68 9493
rect -35 9425 68 9459
rect -35 9391 -7 9425
rect 27 9391 68 9425
rect -35 9357 68 9391
rect -35 9323 -7 9357
rect 27 9323 68 9357
rect -35 9289 68 9323
rect -35 9255 -7 9289
rect 27 9255 68 9289
rect -35 9221 68 9255
rect -35 9187 -7 9221
rect 27 9187 68 9221
rect -35 9153 68 9187
rect -35 9119 -7 9153
rect 27 9119 68 9153
rect -35 9085 68 9119
rect -35 9051 -7 9085
rect 27 9051 68 9085
rect -35 9017 68 9051
rect -35 8983 -7 9017
rect 27 8983 68 9017
rect -35 8949 68 8983
rect -35 8915 -7 8949
rect 27 8915 68 8949
rect -35 8881 68 8915
rect -35 8847 -7 8881
rect 27 8847 68 8881
rect -35 8813 68 8847
rect -35 8779 -7 8813
rect 27 8779 68 8813
rect -35 8745 68 8779
rect -35 8711 -7 8745
rect 27 8711 68 8745
rect -35 8677 68 8711
rect -35 8643 -7 8677
rect 27 8643 68 8677
rect -35 8609 68 8643
rect -35 8575 -7 8609
rect 27 8575 68 8609
rect -35 8541 68 8575
rect -35 8507 -7 8541
rect 27 8507 68 8541
rect -35 8473 68 8507
rect -35 8439 -7 8473
rect 27 8439 68 8473
rect -35 8405 68 8439
rect -35 8371 -7 8405
rect 27 8371 68 8405
rect -35 8337 68 8371
rect -35 8303 -7 8337
rect 27 8303 68 8337
rect -35 8269 68 8303
rect -35 8235 -7 8269
rect 27 8235 68 8269
rect -35 8201 68 8235
rect -35 8167 -7 8201
rect 27 8167 68 8201
rect -35 8133 68 8167
rect -35 8099 -7 8133
rect 27 8099 68 8133
rect -35 8065 68 8099
rect -35 8031 -7 8065
rect 27 8031 68 8065
rect -35 7997 68 8031
rect -35 7963 -7 7997
rect 27 7963 68 7997
rect -35 7929 68 7963
rect -35 7895 -7 7929
rect 27 7895 68 7929
rect -35 7861 68 7895
rect -35 7827 -7 7861
rect 27 7827 68 7861
rect -35 7793 68 7827
rect -35 7759 -7 7793
rect 27 7759 68 7793
rect -35 7725 68 7759
rect -35 7691 -7 7725
rect 27 7691 68 7725
rect -35 7657 68 7691
rect -35 7623 -7 7657
rect 27 7623 68 7657
rect -35 7589 68 7623
rect -35 7555 -7 7589
rect 27 7555 68 7589
rect -35 7521 68 7555
rect -35 7487 -7 7521
rect 27 7487 68 7521
rect -35 7453 68 7487
rect -35 7419 -7 7453
rect 27 7419 68 7453
rect -35 7385 68 7419
rect -35 7351 -7 7385
rect 27 7351 68 7385
rect -35 7317 68 7351
rect -35 7283 -7 7317
rect 27 7283 68 7317
rect -35 7249 68 7283
rect -35 7215 -7 7249
rect 27 7215 68 7249
rect -35 7181 68 7215
rect -35 7147 -7 7181
rect 27 7147 68 7181
rect -35 7113 68 7147
rect -35 7079 -7 7113
rect 27 7079 68 7113
rect -35 7045 68 7079
rect -35 7011 -7 7045
rect 27 7011 68 7045
rect -35 6977 68 7011
rect -35 6943 -7 6977
rect 27 6943 68 6977
rect -35 6909 68 6943
rect -35 6875 -7 6909
rect 27 6875 68 6909
rect -35 6841 68 6875
rect -35 6807 -7 6841
rect 27 6807 68 6841
rect -35 6773 68 6807
rect -35 6739 -7 6773
rect 27 6739 68 6773
rect -35 6705 68 6739
rect -35 6671 -7 6705
rect 27 6671 68 6705
rect -35 6637 68 6671
rect -35 6603 -7 6637
rect 27 6603 68 6637
rect -35 6569 68 6603
rect -35 6535 -7 6569
rect 27 6535 68 6569
rect -35 6501 68 6535
rect -35 6467 -7 6501
rect 27 6467 68 6501
rect -35 6433 68 6467
rect -35 6399 -7 6433
rect 27 6399 68 6433
rect -35 6365 68 6399
rect -35 6331 -7 6365
rect 27 6331 68 6365
rect -35 6297 68 6331
rect -35 6263 -7 6297
rect 27 6263 68 6297
rect -35 6229 68 6263
rect -35 6195 -7 6229
rect 27 6195 68 6229
rect -35 6161 68 6195
rect -35 6127 -7 6161
rect 27 6127 68 6161
rect -35 6093 68 6127
rect -35 6059 -7 6093
rect 27 6059 68 6093
rect -35 6025 68 6059
rect -35 5991 -7 6025
rect 27 5991 68 6025
rect -35 5957 68 5991
rect -35 5923 -7 5957
rect 27 5923 68 5957
rect -35 5889 68 5923
rect -35 5855 -7 5889
rect 27 5855 68 5889
rect -35 5821 68 5855
rect -35 5787 -7 5821
rect 27 5787 68 5821
rect -35 5753 68 5787
rect -35 5719 -7 5753
rect 27 5719 68 5753
rect -35 5685 68 5719
rect -35 5651 -7 5685
rect 27 5651 68 5685
rect -35 5617 68 5651
rect -35 5583 -7 5617
rect 27 5583 68 5617
rect -35 5549 68 5583
rect -35 5515 -7 5549
rect 27 5515 68 5549
rect -35 5481 68 5515
rect -35 5447 -7 5481
rect 27 5447 68 5481
rect -35 5413 68 5447
rect -35 5379 -7 5413
rect 27 5379 68 5413
rect -35 5345 68 5379
rect -35 5311 -7 5345
rect 27 5311 68 5345
rect -35 5277 68 5311
rect -35 5243 -7 5277
rect 27 5243 68 5277
rect -35 5209 68 5243
rect -35 5175 -7 5209
rect 27 5175 68 5209
rect -35 5141 68 5175
rect -35 5107 -7 5141
rect 27 5107 68 5141
rect -35 5073 68 5107
rect -35 5039 -7 5073
rect 27 5039 68 5073
rect -35 5010 68 5039
rect -35 5005 882 5010
rect -35 4971 -7 5005
rect 27 4986 882 5005
rect 27 4971 68 4986
rect -35 4952 68 4971
rect 102 4976 882 4986
rect -35 4937 102 4952
rect -35 4903 -7 4937
rect 27 4918 102 4937
rect 27 4903 68 4918
rect -35 4884 68 4903
rect -35 4869 102 4884
rect -35 4835 -7 4869
rect 27 4850 102 4869
rect 27 4835 68 4850
rect -35 4816 68 4835
rect -35 4801 102 4816
rect -35 4767 -7 4801
rect 27 4782 102 4801
rect 27 4767 68 4782
rect -35 4748 68 4767
rect -35 4733 102 4748
rect -35 4699 -7 4733
rect 27 4714 102 4733
rect 27 4699 68 4714
rect -35 4680 68 4699
rect -35 4665 102 4680
rect -35 4631 -7 4665
rect 27 4646 102 4665
rect 27 4631 68 4646
rect -35 4612 68 4631
rect -35 4597 102 4612
rect -35 4563 -7 4597
rect 27 4578 102 4597
rect 27 4563 68 4578
rect -35 4544 68 4563
rect -35 4529 102 4544
rect -35 4495 -7 4529
rect 27 4510 102 4529
rect 27 4495 68 4510
rect -35 4476 68 4495
rect -35 4461 102 4476
rect -35 4427 -7 4461
rect 27 4442 102 4461
rect 27 4427 68 4442
rect -35 4408 68 4427
rect -35 4393 102 4408
rect -35 4359 -7 4393
rect 27 4374 102 4393
rect 27 4359 68 4374
rect -35 4340 68 4359
rect -35 4325 102 4340
rect -35 4291 -7 4325
rect 27 4306 102 4325
rect 27 4291 68 4306
rect -35 4272 68 4291
rect -35 4257 102 4272
rect -35 4223 -7 4257
rect 27 4238 102 4257
rect 27 4223 68 4238
rect -35 4204 68 4223
rect -35 4189 102 4204
rect -35 4155 -7 4189
rect 27 4170 102 4189
rect 27 4155 68 4170
rect -35 4136 68 4155
rect -35 4121 102 4136
rect -35 4087 -7 4121
rect 27 4102 102 4121
rect 27 4087 68 4102
rect -35 4068 68 4087
rect -35 4053 102 4068
rect -35 4019 -7 4053
rect 27 4034 102 4053
rect 27 4019 68 4034
rect -35 4000 68 4019
rect -35 3985 102 4000
rect -35 3951 -7 3985
rect 27 3966 102 3985
rect 27 3951 68 3966
rect -35 3932 68 3951
rect -35 3917 102 3932
rect -35 3883 -7 3917
rect 27 3898 102 3917
rect 27 3883 68 3898
rect -35 3864 68 3883
rect -35 3849 102 3864
rect -35 3815 -7 3849
rect 27 3830 102 3849
rect 27 3815 68 3830
rect -35 3796 68 3815
rect -35 3781 102 3796
rect -35 3747 -7 3781
rect 27 3762 102 3781
rect 27 3747 68 3762
rect -35 3728 68 3747
rect -35 3713 102 3728
rect -35 3679 -7 3713
rect 27 3694 102 3713
rect 27 3679 68 3694
rect -35 3660 68 3679
rect -35 3645 102 3660
rect -35 3611 -7 3645
rect 27 3626 102 3645
rect 27 3611 68 3626
rect -35 3592 68 3611
rect -35 3577 102 3592
rect -35 3543 -7 3577
rect 27 3558 102 3577
rect 27 3543 68 3558
rect -35 3524 68 3543
rect -35 3508 102 3524
rect -35 3474 -7 3508
rect 27 3490 102 3508
rect 27 3474 68 3490
rect -35 3456 68 3474
rect -35 3439 102 3456
rect -35 3405 -7 3439
rect 27 3422 102 3439
rect 27 3405 68 3422
rect -35 3388 68 3405
rect -35 3370 102 3388
rect -35 3336 -7 3370
rect 27 3354 102 3370
rect 27 3336 68 3354
rect -35 3320 68 3336
rect -35 3301 102 3320
rect -35 3267 -7 3301
rect 27 3286 102 3301
rect 27 3267 68 3286
rect -35 3252 68 3267
rect -35 3232 102 3252
rect -35 3198 -7 3232
rect 27 3218 102 3232
rect 27 3198 68 3218
rect -35 3184 68 3198
rect -35 3163 102 3184
rect -35 3129 -7 3163
rect 27 3150 102 3163
rect 27 3129 68 3150
rect -35 3116 68 3129
rect -35 3094 102 3116
rect -35 3060 -7 3094
rect 27 3082 102 3094
rect 27 3060 68 3082
rect -35 3048 68 3060
rect -35 3025 102 3048
rect -35 2991 -7 3025
rect 27 3014 102 3025
rect 27 2991 68 3014
rect -35 2980 68 2991
rect -35 2956 102 2980
rect -35 2922 -7 2956
rect 27 2946 102 2956
rect 27 2922 68 2946
rect -35 2912 68 2922
rect -35 2887 102 2912
rect -35 2853 -7 2887
rect 27 2878 102 2887
rect 27 2853 68 2878
rect -35 2844 68 2853
rect -35 2818 102 2844
rect -35 2784 -7 2818
rect 27 2810 102 2818
rect 27 2784 68 2810
rect -35 2776 68 2784
rect -35 2749 102 2776
rect -35 2715 -7 2749
rect 27 2742 102 2749
rect 27 2715 68 2742
rect -35 2708 68 2715
rect -35 2680 102 2708
rect -35 2646 -7 2680
rect 27 2674 102 2680
rect 27 2646 68 2674
rect -35 2640 68 2646
rect -35 2611 102 2640
rect -35 2577 -7 2611
rect 27 2606 102 2611
rect 27 2577 68 2606
rect -35 2572 68 2577
rect -35 2542 102 2572
rect -35 2508 -7 2542
rect 27 2538 102 2542
rect 27 2508 68 2538
rect -35 2504 68 2508
rect -35 2473 102 2504
rect -35 2439 -7 2473
rect 27 2470 102 2473
rect 27 2439 68 2470
rect -35 2436 68 2439
rect -35 2404 102 2436
rect -35 2370 -7 2404
rect 27 2402 102 2404
rect 27 2370 68 2402
rect -35 2368 68 2370
rect -35 2335 102 2368
rect -35 2301 -7 2335
rect 27 2334 102 2335
rect 27 2301 68 2334
rect -35 2300 68 2301
rect -35 2266 102 2300
rect -35 2232 -7 2266
rect 27 2232 68 2266
rect -35 2198 102 2232
rect -35 2197 68 2198
rect -35 2163 -7 2197
rect 27 2164 68 2197
rect 27 2163 102 2164
rect -35 2130 102 2163
rect -35 2128 68 2130
rect -35 2094 -7 2128
rect 27 2096 68 2128
rect 27 2094 102 2096
rect -35 2062 102 2094
rect -35 2059 68 2062
rect -35 2025 -7 2059
rect 27 2028 68 2059
rect 27 2025 102 2028
rect -35 1994 102 2025
rect -35 1990 68 1994
rect -35 1956 -7 1990
rect 27 1960 68 1990
rect 27 1956 102 1960
rect -35 1926 102 1956
rect -35 1921 68 1926
rect -35 1887 -7 1921
rect 27 1892 68 1921
rect 27 1887 102 1892
rect -35 1858 102 1887
rect -35 1852 68 1858
rect -35 1818 -7 1852
rect 27 1824 68 1852
rect 27 1818 102 1824
rect -35 1790 102 1818
rect -35 1783 68 1790
rect -35 1749 -7 1783
rect 27 1756 68 1783
rect 27 1749 102 1756
rect -35 1722 102 1749
rect -35 1714 68 1722
rect -35 1680 -7 1714
rect 27 1688 68 1714
rect 27 1680 102 1688
rect -35 1654 102 1680
rect -35 1645 68 1654
rect -35 1611 -7 1645
rect 27 1620 68 1645
rect 27 1611 102 1620
rect -35 1586 102 1611
rect -35 1576 68 1586
rect -35 1542 -7 1576
rect 27 1552 68 1576
rect 27 1542 102 1552
rect -35 1518 102 1542
rect -35 1507 68 1518
rect -35 1473 -7 1507
rect 27 1484 68 1507
rect 27 1473 102 1484
rect -35 1450 102 1473
rect -35 1438 68 1450
rect -35 1404 -7 1438
rect 27 1416 68 1438
rect 27 1404 102 1416
rect -35 1381 102 1404
rect -35 1369 68 1381
rect -35 1335 -7 1369
rect 27 1347 68 1369
rect 27 1335 102 1347
rect -35 1312 102 1335
rect -35 1300 68 1312
rect -35 1266 -7 1300
rect 27 1278 68 1300
rect 27 1266 102 1278
rect -35 1243 102 1266
rect -35 1231 68 1243
rect -35 1197 -7 1231
rect 27 1209 68 1231
rect 27 1197 102 1209
rect -35 1174 102 1197
rect -35 1162 68 1174
rect -35 1128 -7 1162
rect 27 1140 68 1162
rect 27 1128 102 1140
rect -35 1105 102 1128
rect -35 1093 68 1105
rect -35 1059 -7 1093
rect 27 1071 68 1093
rect 27 1059 102 1071
rect -35 1036 102 1059
rect -35 1024 68 1036
rect -35 990 -7 1024
rect 27 1002 68 1024
rect 27 990 102 1002
rect -35 967 102 990
rect -35 955 68 967
rect -35 921 -7 955
rect 27 933 68 955
rect 27 921 102 933
rect -35 898 102 921
rect -35 886 68 898
rect -35 852 -7 886
rect 27 864 68 886
rect 27 852 102 864
rect -35 829 102 852
rect -35 817 68 829
rect -35 783 -7 817
rect 27 795 68 817
rect 27 783 102 795
rect -35 760 102 783
rect -35 748 68 760
rect -35 714 -7 748
rect 27 726 68 748
rect 27 714 102 726
rect -35 691 102 714
rect -35 679 68 691
rect -35 645 -7 679
rect 27 657 68 679
rect 27 645 102 657
rect -35 622 102 645
rect -35 610 68 622
rect -35 576 -7 610
rect 27 588 68 610
rect 27 576 102 588
rect -35 553 102 576
rect -35 541 68 553
rect -35 507 -7 541
rect 27 519 68 541
rect 27 507 102 519
rect -35 484 102 507
rect -35 472 68 484
rect -35 438 -7 472
rect 27 450 68 472
rect 27 438 102 450
rect -35 415 102 438
rect -35 403 68 415
rect -35 369 -7 403
rect 27 381 68 403
rect 27 369 102 381
rect -35 346 102 369
rect -35 334 68 346
rect -35 300 -7 334
rect 27 312 68 334
rect 27 300 102 312
rect -35 277 102 300
rect -35 265 68 277
rect -35 231 -7 265
rect 27 243 68 265
rect 27 231 102 243
rect -35 208 102 231
rect -35 196 68 208
rect -35 162 -7 196
rect 27 174 68 196
rect 27 162 102 174
rect -35 127 102 162
rect -35 93 -7 127
rect 27 102 102 127
rect 848 141 882 4976
rect 848 102 931 141
rect 27 93 92 102
rect -35 68 92 93
rect 126 68 161 102
rect 195 68 230 102
rect 264 68 300 102
rect 334 68 370 102
rect 404 68 440 102
rect 474 68 510 102
rect 544 68 580 102
rect 614 68 650 102
rect 684 68 720 102
rect 754 68 790 102
rect 824 68 931 102
rect -35 58 931 68
rect -35 24 -7 58
rect 27 34 931 58
rect 27 24 92 34
rect -35 0 92 24
rect 126 0 161 34
rect 195 0 230 34
rect 264 0 300 34
rect 334 0 370 34
rect 404 0 440 34
rect 474 0 510 34
rect 544 0 580 34
rect 614 0 650 34
rect 684 0 720 34
rect 754 0 790 34
rect 824 0 931 34
rect -35 -34 931 0
<< mvpsubdiffcont >>
rect 278 4788 312 4822
rect 391 4788 425 4822
rect 525 4788 559 4822
rect 662 4764 696 4798
rect 254 4694 288 4728
rect 254 4625 288 4659
rect 254 4556 288 4590
rect 254 4487 288 4521
rect 254 4418 288 4452
rect 254 4349 288 4383
rect 254 4280 288 4314
rect 254 4211 288 4245
rect 254 4142 288 4176
rect 254 4073 288 4107
rect 254 4004 288 4038
rect 254 3935 288 3969
rect 254 3866 288 3900
rect 254 3797 288 3831
rect 254 3728 288 3762
rect 662 4695 696 4729
rect 662 4626 696 4660
rect 662 4557 696 4591
rect 662 4488 696 4522
rect 662 4419 696 4453
rect 662 4350 696 4384
rect 662 4281 696 4315
rect 662 4212 696 4246
rect 662 4143 696 4177
rect 662 4074 696 4108
rect 662 4005 696 4039
rect 662 3936 696 3970
rect 662 3867 696 3901
rect 662 3798 696 3832
rect 662 3729 696 3763
rect 254 3659 288 3693
rect 254 3590 288 3624
rect 662 3660 696 3694
rect 254 3521 288 3555
rect 254 3452 288 3486
rect 254 3383 288 3417
rect 254 3314 288 3348
rect 254 3245 288 3279
rect 254 3176 288 3210
rect 254 3107 288 3141
rect 254 3038 288 3072
rect 254 2969 288 3003
rect 254 2900 288 2934
rect 254 2831 288 2865
rect 254 2762 288 2796
rect 254 2693 288 2727
rect 254 2624 288 2658
rect 662 3591 696 3625
rect 662 3522 696 3556
rect 662 3453 696 3487
rect 662 3384 696 3418
rect 662 3315 696 3349
rect 662 3246 696 3280
rect 662 3177 696 3211
rect 662 3108 696 3142
rect 662 3039 696 3073
rect 662 2970 696 3004
rect 662 2901 696 2935
rect 662 2832 696 2866
rect 662 2763 696 2797
rect 662 2694 696 2728
rect 662 2625 696 2659
rect 254 2555 288 2589
rect 254 2486 288 2520
rect 662 2556 696 2590
rect 662 2487 696 2521
rect 254 2417 288 2451
rect 254 2348 288 2382
rect 254 2279 288 2313
rect 254 2210 288 2244
rect 254 2141 288 2175
rect 254 2072 288 2106
rect 254 2003 288 2037
rect 254 1934 288 1968
rect 254 1865 288 1899
rect 254 1796 288 1830
rect 254 1727 288 1761
rect 254 1658 288 1692
rect 254 1589 288 1623
rect 254 1520 288 1554
rect 254 1451 288 1485
rect 662 2418 696 2452
rect 662 2349 696 2383
rect 662 2280 696 2314
rect 662 2211 696 2245
rect 662 2142 696 2176
rect 662 2073 696 2107
rect 662 2004 696 2038
rect 662 1935 696 1969
rect 662 1866 696 1900
rect 662 1797 696 1831
rect 662 1728 696 1762
rect 662 1659 696 1693
rect 662 1590 696 1624
rect 662 1521 696 1555
rect 254 1382 288 1416
rect 662 1452 696 1486
rect 662 1383 696 1417
rect 254 1313 288 1347
rect 254 1244 288 1278
rect 254 1175 288 1209
rect 254 1106 288 1140
rect 254 1037 288 1071
rect 254 968 288 1002
rect 254 899 288 933
rect 254 830 288 864
rect 254 761 288 795
rect 254 692 288 726
rect 254 623 288 657
rect 254 554 288 588
rect 254 485 288 519
rect 254 416 288 450
rect 254 347 288 381
rect 662 1314 696 1348
rect 662 1245 696 1279
rect 662 1176 696 1210
rect 662 1107 696 1141
rect 662 1038 696 1072
rect 662 969 696 1003
rect 662 900 696 934
rect 662 831 696 865
rect 662 762 696 796
rect 662 693 696 727
rect 662 624 696 658
rect 662 555 696 589
rect 662 486 696 520
rect 662 417 696 451
rect 662 348 696 382
rect 254 278 288 312
rect 352 254 386 288
rect 423 254 457 288
rect 494 254 528 288
rect 566 254 600 288
rect 638 254 672 288
<< mvnsubdiffcont >>
rect -7 12179 27 12213
rect -7 12111 27 12145
rect -7 12043 27 12077
rect -7 11975 27 12009
rect -7 11907 27 11941
rect -7 11839 27 11873
rect -7 11771 27 11805
rect -7 11703 27 11737
rect -7 11635 27 11669
rect -7 11567 27 11601
rect -7 11499 27 11533
rect -7 11431 27 11465
rect -7 11363 27 11397
rect -7 11295 27 11329
rect -7 11227 27 11261
rect -7 11159 27 11193
rect -7 11091 27 11125
rect -7 11023 27 11057
rect -7 10955 27 10989
rect -7 10887 27 10921
rect -7 10819 27 10853
rect -7 10751 27 10785
rect -7 10683 27 10717
rect -7 10615 27 10649
rect -7 10547 27 10581
rect -7 10479 27 10513
rect -7 10411 27 10445
rect -7 10343 27 10377
rect -7 10275 27 10309
rect -7 10207 27 10241
rect -7 10139 27 10173
rect -7 10071 27 10105
rect -7 10003 27 10037
rect -7 9935 27 9969
rect -7 9867 27 9901
rect -7 9799 27 9833
rect -7 9731 27 9765
rect -7 9663 27 9697
rect -7 9595 27 9629
rect -7 9527 27 9561
rect -7 9459 27 9493
rect -7 9391 27 9425
rect -7 9323 27 9357
rect -7 9255 27 9289
rect -7 9187 27 9221
rect -7 9119 27 9153
rect -7 9051 27 9085
rect -7 8983 27 9017
rect -7 8915 27 8949
rect -7 8847 27 8881
rect -7 8779 27 8813
rect -7 8711 27 8745
rect -7 8643 27 8677
rect -7 8575 27 8609
rect -7 8507 27 8541
rect -7 8439 27 8473
rect -7 8371 27 8405
rect -7 8303 27 8337
rect -7 8235 27 8269
rect -7 8167 27 8201
rect -7 8099 27 8133
rect -7 8031 27 8065
rect -7 7963 27 7997
rect -7 7895 27 7929
rect -7 7827 27 7861
rect -7 7759 27 7793
rect -7 7691 27 7725
rect -7 7623 27 7657
rect -7 7555 27 7589
rect -7 7487 27 7521
rect -7 7419 27 7453
rect -7 7351 27 7385
rect -7 7283 27 7317
rect -7 7215 27 7249
rect -7 7147 27 7181
rect -7 7079 27 7113
rect -7 7011 27 7045
rect -7 6943 27 6977
rect -7 6875 27 6909
rect -7 6807 27 6841
rect -7 6739 27 6773
rect -7 6671 27 6705
rect -7 6603 27 6637
rect -7 6535 27 6569
rect -7 6467 27 6501
rect -7 6399 27 6433
rect -7 6331 27 6365
rect -7 6263 27 6297
rect -7 6195 27 6229
rect -7 6127 27 6161
rect -7 6059 27 6093
rect -7 5991 27 6025
rect -7 5923 27 5957
rect -7 5855 27 5889
rect -7 5787 27 5821
rect -7 5719 27 5753
rect -7 5651 27 5685
rect -7 5583 27 5617
rect -7 5515 27 5549
rect -7 5447 27 5481
rect -7 5379 27 5413
rect -7 5311 27 5345
rect -7 5243 27 5277
rect -7 5175 27 5209
rect -7 5107 27 5141
rect -7 5039 27 5073
rect -7 4971 27 5005
rect 68 4952 102 4986
rect -7 4903 27 4937
rect 68 4884 102 4918
rect -7 4835 27 4869
rect 68 4816 102 4850
rect -7 4767 27 4801
rect 68 4748 102 4782
rect -7 4699 27 4733
rect 68 4680 102 4714
rect -7 4631 27 4665
rect 68 4612 102 4646
rect -7 4563 27 4597
rect 68 4544 102 4578
rect -7 4495 27 4529
rect 68 4476 102 4510
rect -7 4427 27 4461
rect 68 4408 102 4442
rect -7 4359 27 4393
rect 68 4340 102 4374
rect -7 4291 27 4325
rect 68 4272 102 4306
rect -7 4223 27 4257
rect 68 4204 102 4238
rect -7 4155 27 4189
rect 68 4136 102 4170
rect -7 4087 27 4121
rect 68 4068 102 4102
rect -7 4019 27 4053
rect 68 4000 102 4034
rect -7 3951 27 3985
rect 68 3932 102 3966
rect -7 3883 27 3917
rect 68 3864 102 3898
rect -7 3815 27 3849
rect 68 3796 102 3830
rect -7 3747 27 3781
rect 68 3728 102 3762
rect -7 3679 27 3713
rect 68 3660 102 3694
rect -7 3611 27 3645
rect 68 3592 102 3626
rect -7 3543 27 3577
rect 68 3524 102 3558
rect -7 3474 27 3508
rect 68 3456 102 3490
rect -7 3405 27 3439
rect 68 3388 102 3422
rect -7 3336 27 3370
rect 68 3320 102 3354
rect -7 3267 27 3301
rect 68 3252 102 3286
rect -7 3198 27 3232
rect 68 3184 102 3218
rect -7 3129 27 3163
rect 68 3116 102 3150
rect -7 3060 27 3094
rect 68 3048 102 3082
rect -7 2991 27 3025
rect 68 2980 102 3014
rect -7 2922 27 2956
rect 68 2912 102 2946
rect -7 2853 27 2887
rect 68 2844 102 2878
rect -7 2784 27 2818
rect 68 2776 102 2810
rect -7 2715 27 2749
rect 68 2708 102 2742
rect -7 2646 27 2680
rect 68 2640 102 2674
rect -7 2577 27 2611
rect 68 2572 102 2606
rect -7 2508 27 2542
rect 68 2504 102 2538
rect -7 2439 27 2473
rect 68 2436 102 2470
rect -7 2370 27 2404
rect 68 2368 102 2402
rect -7 2301 27 2335
rect 68 2300 102 2334
rect -7 2232 27 2266
rect 68 2232 102 2266
rect -7 2163 27 2197
rect 68 2164 102 2198
rect -7 2094 27 2128
rect 68 2096 102 2130
rect -7 2025 27 2059
rect 68 2028 102 2062
rect -7 1956 27 1990
rect 68 1960 102 1994
rect -7 1887 27 1921
rect 68 1892 102 1926
rect -7 1818 27 1852
rect 68 1824 102 1858
rect -7 1749 27 1783
rect 68 1756 102 1790
rect -7 1680 27 1714
rect 68 1688 102 1722
rect -7 1611 27 1645
rect 68 1620 102 1654
rect -7 1542 27 1576
rect 68 1552 102 1586
rect -7 1473 27 1507
rect 68 1484 102 1518
rect -7 1404 27 1438
rect 68 1416 102 1450
rect -7 1335 27 1369
rect 68 1347 102 1381
rect -7 1266 27 1300
rect 68 1278 102 1312
rect -7 1197 27 1231
rect 68 1209 102 1243
rect -7 1128 27 1162
rect 68 1140 102 1174
rect -7 1059 27 1093
rect 68 1071 102 1105
rect -7 990 27 1024
rect 68 1002 102 1036
rect -7 921 27 955
rect 68 933 102 967
rect -7 852 27 886
rect 68 864 102 898
rect -7 783 27 817
rect 68 795 102 829
rect -7 714 27 748
rect 68 726 102 760
rect -7 645 27 679
rect 68 657 102 691
rect -7 576 27 610
rect 68 588 102 622
rect -7 507 27 541
rect 68 519 102 553
rect -7 438 27 472
rect 68 450 102 484
rect -7 369 27 403
rect 68 381 102 415
rect -7 300 27 334
rect 68 312 102 346
rect -7 231 27 265
rect 68 243 102 277
rect -7 162 27 196
rect 68 174 102 208
rect -7 93 27 127
rect 92 68 126 102
rect 161 68 195 102
rect 230 68 264 102
rect 300 68 334 102
rect 370 68 404 102
rect 440 68 474 102
rect 510 68 544 102
rect 580 68 614 102
rect 650 68 684 102
rect 720 68 754 102
rect 790 68 824 102
rect -7 24 27 58
rect 92 0 126 34
rect 161 0 195 34
rect 230 0 264 34
rect 300 0 334 34
rect 370 0 404 34
rect 440 0 474 34
rect 510 0 544 34
rect 580 0 614 34
rect 650 0 684 34
rect 720 0 754 34
rect 790 0 824 34
<< poly >>
rect 415 4714 535 4740
rect 415 3674 535 3714
rect 415 3640 472 3674
rect 506 3640 535 3674
rect 415 3593 535 3640
rect 415 2553 535 2593
rect 415 2519 472 2553
rect 506 2519 535 2553
rect 415 2472 535 2519
rect 415 1434 535 1472
rect 415 1400 472 1434
rect 506 1400 535 1434
rect 415 1362 535 1400
rect 415 336 535 362
<< polycont >>
rect 472 3640 506 3674
rect 472 2519 506 2553
rect 472 1400 506 1434
<< locali >>
rect -35 12213 55 12237
rect -35 12179 -7 12213
rect 27 12179 55 12213
rect -35 12145 55 12179
rect -35 12129 -7 12145
rect 27 12129 55 12145
rect -35 12095 -20 12129
rect 27 12111 52 12129
rect 14 12095 52 12111
rect -35 12077 86 12095
rect -35 12055 -7 12077
rect 27 12055 86 12077
rect -35 12021 -20 12055
rect 27 12043 52 12055
rect 14 12021 52 12043
rect -35 12009 86 12021
rect 197 12010 246 12044
rect 280 12010 329 12044
rect 363 12010 412 12044
rect 446 12010 496 12044
rect 530 12010 580 12044
rect 614 12010 664 12044
rect 698 12010 770 12044
rect -35 11981 -7 12009
rect 27 11981 86 12009
rect -35 11947 -20 11981
rect 27 11975 52 11981
rect 14 11947 52 11975
rect 736 11972 770 12010
rect -35 11941 86 11947
rect -35 11907 -7 11941
rect 27 11907 86 11941
rect -35 11873 -20 11907
rect 14 11873 52 11907
rect -35 11839 -7 11873
rect 27 11839 86 11873
rect -35 11833 86 11839
rect -35 11799 -20 11833
rect 14 11805 52 11833
rect 27 11799 52 11805
rect -35 11771 -7 11799
rect 27 11771 86 11799
rect -35 11759 86 11771
rect -35 11725 -20 11759
rect 14 11737 52 11759
rect 27 11725 52 11737
rect -35 11703 -7 11725
rect 27 11703 86 11725
rect -35 11685 86 11703
rect -35 11651 -20 11685
rect 14 11669 52 11685
rect 27 11651 52 11669
rect -35 11635 -7 11651
rect 27 11635 86 11651
rect -35 11611 86 11635
rect -35 11577 -20 11611
rect 14 11601 52 11611
rect 27 11577 52 11601
rect -35 11567 -7 11577
rect 27 11567 86 11577
rect -35 11537 86 11567
rect -35 11503 -20 11537
rect 14 11533 52 11537
rect 27 11503 52 11533
rect -35 11499 -7 11503
rect 27 11499 86 11503
rect -35 11465 86 11499
rect -35 11463 -7 11465
rect 27 11463 86 11465
rect -35 11429 -20 11463
rect 27 11431 52 11463
rect 14 11429 52 11431
rect -35 11397 86 11429
rect -35 11389 -7 11397
rect 27 11389 86 11397
rect -35 11355 -20 11389
rect 27 11363 52 11389
rect 14 11355 52 11363
rect -35 11329 86 11355
rect -35 11315 -7 11329
rect 27 11315 86 11329
rect -35 11281 -20 11315
rect 27 11295 52 11315
rect 14 11281 52 11295
rect -35 11261 86 11281
rect -35 11241 -7 11261
rect 27 11241 86 11261
rect -35 11207 -20 11241
rect 27 11227 52 11241
rect 14 11207 52 11227
rect -35 11193 86 11207
rect -35 11167 -7 11193
rect 27 11167 86 11193
rect -35 11133 -20 11167
rect 27 11159 52 11167
rect 14 11133 52 11159
rect -35 11125 86 11133
rect -35 11093 -7 11125
rect 27 11093 86 11125
rect -35 11059 -20 11093
rect 27 11091 52 11093
rect 14 11059 52 11091
rect -35 11057 86 11059
rect -35 11023 -7 11057
rect 27 11023 86 11057
rect -35 11019 86 11023
rect -35 10985 -20 11019
rect 14 10989 52 11019
rect 27 10985 52 10989
rect -35 10955 -7 10985
rect 27 10955 86 10985
rect -35 10945 86 10955
rect -35 10911 -20 10945
rect 14 10921 52 10945
rect 27 10911 52 10921
rect -35 10887 -7 10911
rect 27 10887 86 10911
rect -35 10871 86 10887
rect -35 10837 -20 10871
rect 14 10853 52 10871
rect 27 10837 52 10853
rect -35 10819 -7 10837
rect 27 10819 86 10837
rect -35 10797 86 10819
rect -35 10763 -20 10797
rect 14 10785 52 10797
rect 27 10763 52 10785
rect -35 10751 -7 10763
rect 27 10751 86 10763
rect -35 10723 86 10751
rect -35 10689 -20 10723
rect 14 10717 52 10723
rect 27 10689 52 10717
rect -35 10683 -7 10689
rect 27 10683 86 10689
rect -35 10649 86 10683
rect -35 10615 -20 10649
rect 27 10615 52 10649
rect -35 10581 86 10615
rect -35 10575 -7 10581
rect 27 10575 86 10581
rect -35 10541 -20 10575
rect 27 10547 52 10575
rect 14 10541 52 10547
rect -35 10513 86 10541
rect -35 10502 -7 10513
rect 27 10502 86 10513
rect -35 10468 -20 10502
rect 27 10479 52 10502
rect 14 10468 52 10479
rect 158 11925 230 11959
rect 264 11925 302 11959
rect 336 11925 374 11959
rect 408 11925 446 11959
rect 480 11925 518 11959
rect 552 11925 590 11959
rect 624 11925 696 11959
rect 158 11887 192 11925
rect 158 11811 192 11853
rect 158 11735 192 11777
rect 158 11659 192 11701
rect 158 11583 192 11625
rect 158 11507 192 11549
rect 158 11431 192 11473
rect 158 11355 192 11397
rect 158 11279 192 11321
rect 158 11203 192 11245
rect 158 11127 192 11169
rect 158 11051 192 11093
rect 158 10975 192 11017
rect 158 10899 192 10941
rect 158 10823 192 10865
rect 158 10747 192 10789
rect 158 10672 192 10713
rect 158 10597 192 10638
rect 158 10522 192 10563
rect 662 11887 696 11925
rect 662 11815 696 11853
rect 662 11743 696 11781
rect 662 11671 696 11709
rect 662 11599 696 11637
rect 662 11527 696 11565
rect 662 11455 696 11493
rect 662 11383 696 11421
rect 662 11311 696 11349
rect 662 11239 696 11277
rect 662 11167 696 11205
rect 662 11095 696 11133
rect 662 11023 696 11061
rect 662 10951 696 10989
rect 662 10879 696 10917
rect 662 10807 696 10845
rect 662 10735 696 10773
rect 662 10663 696 10701
rect 662 10591 696 10629
rect 662 10519 696 10557
rect -35 10445 86 10468
rect -35 10429 -7 10445
rect 27 10429 86 10445
rect 662 10447 696 10485
rect -35 10395 -20 10429
rect 27 10411 52 10429
rect 14 10395 52 10411
rect -35 10377 86 10395
rect -35 10356 -7 10377
rect 27 10356 86 10377
rect -35 10322 -20 10356
rect 27 10343 52 10356
rect 14 10322 52 10343
rect -35 10309 86 10322
rect -35 10283 -7 10309
rect 27 10283 86 10309
rect -35 10249 -20 10283
rect 27 10275 52 10283
rect 14 10249 52 10275
rect -35 10241 86 10249
rect -35 10210 -7 10241
rect 27 10210 86 10241
rect -35 10176 -20 10210
rect 27 10207 52 10210
rect 14 10176 52 10207
rect -35 10173 86 10176
rect -35 10139 -7 10173
rect 27 10139 86 10173
rect -35 10137 86 10139
rect -35 10103 -20 10137
rect 14 10105 52 10137
rect 27 10103 52 10105
rect -35 10071 -7 10103
rect 27 10071 86 10103
rect -35 10064 86 10071
rect -35 10030 -20 10064
rect 14 10037 52 10064
rect 27 10030 52 10037
rect -35 10003 -7 10030
rect 27 10003 86 10030
rect -35 9991 86 10003
rect -35 9957 -20 9991
rect 14 9969 52 9991
rect 27 9957 52 9969
rect -35 9935 -7 9957
rect 27 9935 86 9957
rect -35 9918 86 9935
rect -35 9884 -20 9918
rect 14 9901 52 9918
rect 27 9884 52 9901
rect -35 9867 -7 9884
rect 27 9867 86 9884
rect -35 9845 86 9867
rect 192 10405 278 10439
rect 158 10360 312 10405
rect 192 10326 278 10360
rect 158 10281 312 10326
rect 192 10247 278 10281
rect 158 10202 312 10247
rect 192 10168 278 10202
rect 158 10123 312 10168
rect 192 10089 278 10123
rect 158 10043 312 10089
rect 192 10009 278 10043
rect 158 9963 312 10009
rect 192 9929 278 9963
rect 158 9883 312 9929
rect 192 9849 278 9883
rect 662 10375 696 10413
rect 662 10303 696 10341
rect 662 10231 696 10269
rect 662 10159 696 10197
rect 662 10087 696 10125
rect 662 10015 696 10053
rect 662 9943 696 9981
rect 662 9871 696 9909
rect -35 9811 -20 9845
rect 14 9833 52 9845
rect 27 9811 52 9833
rect -35 9799 -7 9811
rect 27 9799 86 9811
rect -35 9772 86 9799
rect -35 9738 -20 9772
rect 14 9765 52 9772
rect 27 9738 52 9765
rect -35 9731 -7 9738
rect 27 9731 86 9738
rect -35 9699 86 9731
rect -35 9665 -20 9699
rect 14 9697 52 9699
rect 27 9665 52 9697
rect -35 9663 -7 9665
rect 27 9663 86 9665
rect -35 9629 86 9663
rect -35 9626 -7 9629
rect 27 9626 86 9629
rect -35 9592 -20 9626
rect 27 9595 52 9626
rect 14 9592 52 9595
rect -35 9561 86 9592
rect -35 9553 -7 9561
rect 27 9553 86 9561
rect -35 9519 -20 9553
rect 27 9527 52 9553
rect 14 9519 52 9527
rect -35 9493 86 9519
rect -35 9480 -7 9493
rect 27 9480 86 9493
rect -35 9446 -20 9480
rect 27 9459 52 9480
rect 14 9446 52 9459
rect 662 9799 696 9837
rect 662 9727 696 9765
rect 662 9655 696 9693
rect 662 9583 696 9621
rect 662 9511 696 9549
rect -35 9425 55 9446
rect -35 9391 -7 9425
rect 27 9391 55 9425
rect -35 9357 55 9391
rect -35 9323 -7 9357
rect 27 9323 55 9357
rect -35 9289 55 9323
rect -35 9255 -7 9289
rect 27 9255 55 9289
rect -35 9221 55 9255
rect -35 9187 -7 9221
rect 27 9187 55 9221
rect -35 9163 55 9187
rect 662 9439 696 9477
rect 662 9367 696 9405
rect 662 9294 696 9333
rect 662 9221 696 9260
rect -35 9129 -20 9163
rect 14 9153 52 9163
rect 27 9129 52 9153
rect -35 9119 -7 9129
rect 27 9119 86 9129
rect -35 9088 86 9119
rect -35 9054 -20 9088
rect 14 9085 52 9088
rect 27 9054 52 9085
rect -35 9051 -7 9054
rect 27 9051 86 9054
rect -35 9017 86 9051
rect -35 9013 -7 9017
rect 27 9013 86 9017
rect -35 8979 -20 9013
rect 27 8983 52 9013
rect 14 8979 52 8983
rect -35 8949 86 8979
rect -35 8938 -7 8949
rect 27 8938 86 8949
rect -35 8904 -20 8938
rect 27 8915 52 8938
rect 14 8904 52 8915
rect -35 8881 86 8904
rect -35 8863 -7 8881
rect 27 8863 86 8881
rect -35 8829 -20 8863
rect 27 8847 52 8863
rect 14 8829 52 8847
rect -35 8813 86 8829
rect -35 8788 -7 8813
rect 27 8788 86 8813
rect -35 8754 -20 8788
rect 27 8779 52 8788
rect 14 8754 52 8779
rect -35 8745 86 8754
rect -35 8713 -7 8745
rect 27 8713 86 8745
rect -35 8679 -20 8713
rect 27 8711 52 8713
rect 14 8679 52 8711
rect -35 8677 86 8679
rect -35 8643 -7 8677
rect 27 8643 86 8677
rect -35 8638 86 8643
rect -35 8604 -20 8638
rect 14 8609 52 8638
rect 27 8604 52 8609
rect 662 9148 696 9187
rect 662 9075 696 9114
rect 662 9002 696 9041
rect 662 8929 696 8968
rect 662 8856 696 8895
rect 662 8783 696 8822
rect 662 8710 696 8749
rect 662 8637 696 8676
rect -35 8575 -7 8604
rect 27 8575 86 8604
rect -35 8563 86 8575
rect -35 8529 -20 8563
rect 14 8541 52 8563
rect 27 8529 52 8541
rect -35 8507 -7 8529
rect 27 8507 86 8529
rect -35 8488 86 8507
rect -35 8454 -20 8488
rect 14 8473 52 8488
rect 27 8454 52 8473
rect -35 8439 -7 8454
rect 27 8439 86 8454
rect -35 8413 86 8439
rect -35 8379 -20 8413
rect 14 8405 52 8413
rect 27 8379 52 8405
rect -35 8371 -7 8379
rect 27 8371 86 8379
rect -35 8338 86 8371
rect -35 8304 -20 8338
rect 14 8337 52 8338
rect 27 8304 52 8337
rect -35 8303 -7 8304
rect 27 8303 86 8304
rect -35 8269 86 8303
rect -35 8263 -7 8269
rect 27 8263 86 8269
rect -35 8229 -20 8263
rect 27 8235 52 8263
rect 14 8229 52 8235
rect -35 8201 86 8229
rect -35 8188 -7 8201
rect 27 8188 86 8201
rect -35 8154 -20 8188
rect 27 8167 52 8188
rect 14 8154 52 8167
rect -35 8133 86 8154
rect -35 8113 -7 8133
rect 27 8113 86 8133
rect -35 8079 -20 8113
rect 27 8099 52 8113
rect 14 8079 52 8099
rect -35 8065 86 8079
rect -35 8038 -7 8065
rect 27 8038 86 8065
rect -35 8004 -20 8038
rect 27 8031 52 8038
rect 14 8004 52 8031
rect 192 8587 278 8621
rect 158 8542 312 8587
rect 192 8508 278 8542
rect 158 8463 312 8508
rect 192 8429 278 8463
rect 158 8384 312 8429
rect 192 8350 278 8384
rect 158 8305 312 8350
rect 192 8271 278 8305
rect 158 8225 312 8271
rect 192 8191 278 8225
rect 158 8145 312 8191
rect 192 8111 278 8145
rect 158 8065 312 8111
rect 192 8031 278 8065
rect 662 8564 696 8603
rect 662 8491 696 8530
rect 662 8418 696 8457
rect 662 8345 696 8384
rect 662 8272 696 8311
rect 662 8199 696 8238
rect 662 8126 696 8165
rect 662 8053 696 8092
rect -35 7997 86 8004
rect -35 7963 -7 7997
rect 27 7963 86 7997
rect -35 7929 -20 7963
rect 14 7929 52 7963
rect -35 7895 -7 7929
rect 27 7895 86 7929
rect -35 7889 86 7895
rect -35 7855 -20 7889
rect 14 7861 52 7889
rect 27 7855 52 7861
rect -35 7827 -7 7855
rect 27 7827 86 7855
rect -35 7815 86 7827
rect -35 7781 -20 7815
rect 14 7793 52 7815
rect 27 7781 52 7793
rect -35 7759 -7 7781
rect 27 7759 86 7781
rect -35 7741 86 7759
rect -35 7707 -20 7741
rect 14 7725 52 7741
rect 27 7707 52 7725
rect -35 7691 -7 7707
rect 27 7691 86 7707
rect -35 7667 86 7691
rect -35 7633 -20 7667
rect 14 7657 52 7667
rect 27 7633 52 7657
rect -35 7623 -7 7633
rect 27 7623 86 7633
rect -35 7593 86 7623
rect -35 7559 -20 7593
rect 14 7589 52 7593
rect 27 7559 52 7589
rect 662 7980 696 8019
rect 662 7907 696 7946
rect 662 7834 696 7873
rect 662 7761 696 7800
rect 662 7688 696 7727
rect 662 7615 696 7654
rect -35 7555 -7 7559
rect 27 7555 55 7559
rect -35 7521 55 7555
rect -35 7487 -7 7521
rect 27 7487 55 7521
rect -35 7453 55 7487
rect -35 7419 -7 7453
rect 27 7419 55 7453
rect -35 7385 55 7419
rect -35 7351 -7 7385
rect 27 7351 55 7385
rect -35 7317 55 7351
rect -35 7283 -7 7317
rect 27 7283 55 7317
rect -35 7268 55 7283
rect 662 7542 696 7581
rect 662 7469 696 7508
rect 662 7396 696 7435
rect 662 7323 696 7362
rect -35 7234 -20 7268
rect 14 7249 52 7268
rect 27 7234 52 7249
rect -35 7215 -7 7234
rect 27 7215 86 7234
rect -35 7194 86 7215
rect -35 7160 -20 7194
rect 14 7181 52 7194
rect 27 7160 52 7181
rect -35 7147 -7 7160
rect 27 7147 86 7160
rect -35 7120 86 7147
rect -35 7086 -20 7120
rect 14 7113 52 7120
rect 27 7086 52 7113
rect -35 7079 -7 7086
rect 27 7079 86 7086
rect -35 7046 86 7079
rect -35 7012 -20 7046
rect 14 7045 52 7046
rect 27 7012 52 7045
rect -35 7011 -7 7012
rect 27 7011 86 7012
rect -35 6977 86 7011
rect -35 6972 -7 6977
rect 27 6972 86 6977
rect -35 6938 -20 6972
rect 27 6943 52 6972
rect 14 6938 52 6943
rect -35 6909 86 6938
rect -35 6898 -7 6909
rect 27 6898 86 6909
rect -35 6864 -20 6898
rect 27 6875 52 6898
rect 14 6864 52 6875
rect -35 6841 86 6864
rect -35 6824 -7 6841
rect 27 6824 86 6841
rect -35 6790 -20 6824
rect 27 6807 52 6824
rect 14 6790 52 6807
rect -35 6773 86 6790
rect -35 6750 -7 6773
rect 27 6750 86 6773
rect -35 6716 -20 6750
rect 27 6739 52 6750
rect 14 6716 52 6739
rect -35 6705 86 6716
rect -35 6676 -7 6705
rect 27 6676 86 6705
rect -35 6642 -20 6676
rect 27 6671 52 6676
rect 14 6642 52 6671
rect -35 6637 86 6642
rect -35 6603 -7 6637
rect 27 6603 86 6637
rect -35 6602 86 6603
rect -35 6568 -20 6602
rect 14 6569 52 6602
rect 27 6568 52 6569
rect -35 6535 -7 6568
rect 27 6535 86 6568
rect -35 6528 86 6535
rect -35 6494 -20 6528
rect 14 6501 52 6528
rect 27 6494 52 6501
rect -35 6467 -7 6494
rect 27 6467 86 6494
rect -35 6454 86 6467
rect -35 6420 -20 6454
rect 14 6433 52 6454
rect 27 6420 52 6433
rect -35 6399 -7 6420
rect 27 6399 86 6420
rect -35 6380 86 6399
rect -35 6346 -20 6380
rect 14 6365 52 6380
rect 27 6346 52 6365
rect -35 6331 -7 6346
rect 27 6331 86 6346
rect -35 6306 86 6331
rect -35 6272 -20 6306
rect 14 6297 52 6306
rect 27 6272 52 6297
rect -35 6263 -7 6272
rect 27 6263 86 6272
rect -35 6233 86 6263
rect -35 6199 -20 6233
rect 14 6229 52 6233
rect 27 6199 52 6229
rect -35 6195 -7 6199
rect 27 6195 86 6199
rect -35 6161 86 6195
rect -35 6160 -7 6161
rect 27 6160 86 6161
rect -35 6126 -20 6160
rect 27 6127 52 6160
rect 14 6126 52 6127
rect -35 6093 86 6126
rect -35 6087 -7 6093
rect 27 6087 86 6093
rect -35 6053 -20 6087
rect 27 6059 52 6087
rect 14 6053 52 6059
rect -35 6025 86 6053
rect -35 6014 -7 6025
rect 27 6014 86 6025
rect -35 5980 -20 6014
rect 27 5991 52 6014
rect 14 5980 52 5991
rect -35 5957 86 5980
rect -35 5941 -7 5957
rect 27 5941 86 5957
rect -35 5907 -20 5941
rect 27 5923 52 5941
rect 14 5907 52 5923
rect -35 5889 86 5907
rect -35 5868 -7 5889
rect 27 5868 86 5889
rect -35 5834 -20 5868
rect 27 5855 52 5868
rect 14 5834 52 5855
rect -35 5821 86 5834
rect -35 5795 -7 5821
rect 27 5795 86 5821
rect -35 5761 -20 5795
rect 27 5787 52 5795
rect 14 5761 52 5787
rect -35 5753 86 5761
rect -35 5722 -7 5753
rect 27 5722 86 5753
rect -35 5688 -20 5722
rect 27 5719 52 5722
rect 14 5688 52 5719
rect -35 5685 86 5688
rect -35 5651 -7 5685
rect 27 5651 86 5685
rect -35 5649 86 5651
rect -35 5615 -20 5649
rect 14 5617 52 5649
rect 27 5615 52 5617
rect -35 5583 -7 5615
rect 27 5583 86 5615
rect -35 5576 86 5583
rect -35 5542 -20 5576
rect 14 5549 52 5576
rect 27 5542 52 5549
rect -35 5515 -7 5542
rect 27 5515 86 5542
rect -35 5503 86 5515
rect -35 5469 -20 5503
rect 14 5481 52 5503
rect 27 5469 52 5481
rect -35 5447 -7 5469
rect 27 5447 86 5469
rect -35 5430 86 5447
rect -35 5396 -20 5430
rect 14 5413 52 5430
rect 27 5396 52 5413
rect -35 5379 -7 5396
rect 27 5379 86 5396
rect -35 5357 86 5379
rect -35 5323 -20 5357
rect 14 5345 52 5357
rect 27 5323 52 5345
rect -35 5311 -7 5323
rect 27 5311 86 5323
rect -35 5284 86 5311
rect -35 5250 -20 5284
rect 14 5277 52 5284
rect 27 5250 52 5277
rect -35 5243 -7 5250
rect 27 5243 86 5250
rect -35 5211 86 5243
rect -35 5177 -20 5211
rect 14 5209 52 5211
rect 27 5177 52 5209
rect -35 5175 -7 5177
rect 27 5175 86 5177
rect -35 5141 86 5175
rect -35 5138 -7 5141
rect 27 5138 86 5141
rect -35 5104 -20 5138
rect 27 5107 52 5138
rect 14 5104 52 5107
rect 159 7239 171 7273
rect 205 7239 217 7273
rect 159 7199 217 7239
rect 159 7165 171 7199
rect 205 7165 217 7199
rect 159 7125 217 7165
rect 159 7091 171 7125
rect 205 7091 217 7125
rect 159 7052 217 7091
rect 159 7018 171 7052
rect 205 7018 217 7052
rect 159 6979 217 7018
rect 159 6945 171 6979
rect 205 6945 217 6979
rect 159 6906 217 6945
rect 159 6872 171 6906
rect 205 6872 217 6906
rect 159 6833 217 6872
rect 159 6799 171 6833
rect 205 6799 217 6833
rect 159 6760 217 6799
rect 159 6726 171 6760
rect 205 6726 217 6760
rect 159 6687 217 6726
rect 159 6653 171 6687
rect 205 6653 217 6687
rect 159 6614 217 6653
rect 159 6580 171 6614
rect 205 6580 217 6614
rect 159 6541 217 6580
rect 159 6507 171 6541
rect 205 6507 217 6541
rect 159 6468 217 6507
rect 159 6434 171 6468
rect 205 6434 217 6468
rect 159 6395 217 6434
rect 159 6361 171 6395
rect 205 6361 217 6395
rect 159 6322 217 6361
rect 159 6288 171 6322
rect 205 6288 217 6322
rect 159 6249 217 6288
rect 159 6215 171 6249
rect 205 6215 217 6249
rect 159 6176 217 6215
rect 159 6142 171 6176
rect 205 6142 217 6176
rect 159 6103 217 6142
rect 159 6069 171 6103
rect 205 6069 217 6103
rect 159 6030 217 6069
rect 159 5996 171 6030
rect 205 5996 217 6030
rect 159 5957 217 5996
rect 159 5923 171 5957
rect 205 5923 217 5957
rect 159 5884 217 5923
rect 159 5850 171 5884
rect 205 5850 217 5884
rect 159 5811 217 5850
rect 159 5777 171 5811
rect 205 5777 217 5811
rect 159 5738 217 5777
rect 159 5704 171 5738
rect 205 5704 217 5738
rect 159 5665 217 5704
rect 159 5631 171 5665
rect 205 5631 217 5665
rect 159 5592 217 5631
rect 159 5558 171 5592
rect 205 5558 217 5592
rect 159 5519 217 5558
rect 159 5485 171 5519
rect 205 5485 217 5519
rect 159 5446 217 5485
rect 159 5412 171 5446
rect 205 5412 217 5446
rect 159 5373 217 5412
rect 159 5339 171 5373
rect 205 5339 217 5373
rect 159 5300 217 5339
rect 159 5266 171 5300
rect 205 5266 217 5300
rect 159 5227 217 5266
rect 159 5193 171 5227
rect 205 5193 217 5227
rect 662 7250 696 7289
rect 662 7177 696 7216
rect 662 7104 696 7143
rect 662 7031 696 7070
rect 662 6958 696 6997
rect 662 6885 696 6924
rect 662 6812 696 6851
rect 662 6739 696 6778
rect 662 6666 696 6705
rect 662 6593 696 6632
rect 662 6520 696 6559
rect 662 6447 696 6486
rect 662 6374 696 6413
rect 662 6301 696 6340
rect 662 6228 696 6267
rect 662 6155 696 6194
rect 662 6082 696 6121
rect 662 6009 696 6048
rect 662 5936 696 5975
rect 662 5863 696 5902
rect 662 5790 696 5829
rect 662 5717 696 5756
rect 662 5644 696 5683
rect 662 5571 696 5610
rect 662 5498 696 5537
rect 662 5425 696 5464
rect 662 5352 696 5391
rect 662 5279 696 5318
rect 662 5207 696 5245
rect 159 5154 217 5193
rect 331 5173 370 5207
rect 404 5173 443 5207
rect 477 5173 516 5207
rect 550 5173 589 5207
rect 623 5173 696 5207
rect 736 11900 770 11938
rect 736 11828 770 11866
rect 736 11756 770 11794
rect 736 11684 770 11722
rect 736 11612 770 11650
rect 736 11540 770 11578
rect 736 11468 770 11506
rect 736 11396 770 11434
rect 736 11324 770 11362
rect 736 11252 770 11290
rect 736 11180 770 11218
rect 736 11108 770 11146
rect 736 11036 770 11074
rect 736 10964 770 11002
rect 736 10892 770 10930
rect 736 10820 770 10858
rect 736 10748 770 10786
rect 736 10676 770 10714
rect 736 10604 770 10642
rect 736 10532 770 10570
rect 736 10460 770 10498
rect 736 10388 770 10426
rect 736 10316 770 10354
rect 736 10244 770 10282
rect 736 10172 770 10210
rect 736 10100 770 10138
rect 736 10028 770 10066
rect 736 9956 770 9994
rect 736 9884 770 9922
rect 736 9812 770 9850
rect 736 9740 770 9778
rect 736 9668 770 9706
rect 736 9596 770 9634
rect 736 9524 770 9562
rect 736 9452 770 9490
rect 736 9380 770 9418
rect 736 9308 770 9346
rect 736 9236 770 9274
rect 736 9164 770 9202
rect 736 9092 770 9130
rect 736 9020 770 9058
rect 736 8948 770 8986
rect 736 8876 770 8914
rect 736 8804 770 8842
rect 736 8732 770 8770
rect 736 8660 770 8698
rect 736 8588 770 8626
rect 736 8516 770 8554
rect 736 8444 770 8482
rect 736 8372 770 8410
rect 736 8300 770 8338
rect 736 8228 770 8266
rect 736 8156 770 8194
rect 736 8084 770 8122
rect 736 8012 770 8050
rect 736 7940 770 7978
rect 736 7868 770 7906
rect 736 7796 770 7834
rect 736 7724 770 7762
rect 736 7652 770 7690
rect 736 7580 770 7618
rect 736 7508 770 7546
rect 736 7436 770 7474
rect 736 7364 770 7402
rect 736 7292 770 7330
rect 736 7220 770 7258
rect 736 7148 770 7186
rect 736 7076 770 7114
rect 736 7004 770 7042
rect 736 6932 770 6970
rect 736 6860 770 6898
rect 736 6788 770 6826
rect 736 6716 770 6754
rect 736 6644 770 6682
rect 736 6572 770 6610
rect 736 6500 770 6538
rect 736 6428 770 6466
rect 736 6356 770 6394
rect 736 6284 770 6322
rect 736 6212 770 6250
rect 736 6140 770 6178
rect 736 6068 770 6106
rect 736 5996 770 6034
rect 736 5924 770 5962
rect 736 5852 770 5890
rect 736 5780 770 5818
rect 736 5708 770 5746
rect 736 5636 770 5674
rect 736 5564 770 5602
rect 736 5492 770 5530
rect 736 5420 770 5458
rect 736 5348 770 5386
rect 736 5275 770 5314
rect 736 5202 770 5241
rect 159 5120 171 5154
rect 205 5120 217 5154
rect 736 5130 770 5168
rect -35 5073 86 5104
rect 331 5096 371 5130
rect 405 5096 444 5130
rect 478 5096 517 5130
rect 551 5096 590 5130
rect 624 5096 663 5130
rect 697 5096 770 5130
rect -35 5065 -7 5073
rect 27 5065 86 5073
rect -35 5031 -20 5065
rect 27 5039 52 5065
rect 14 5031 52 5039
rect -35 5010 86 5031
rect 848 5010 930 12162
rect -44 5005 129 5010
rect -44 4992 -7 5005
rect 27 4992 129 5005
rect -44 4958 -20 4992
rect 27 4971 52 4992
rect 86 4986 129 4992
rect 14 4958 52 4971
rect 102 4976 129 4986
rect 163 4976 205 5010
rect 239 4976 281 5010
rect 315 4976 357 5010
rect 391 4976 433 5010
rect 467 4976 508 5010
rect 542 4976 583 5010
rect 617 4976 658 5010
rect 692 4976 733 5010
rect 767 4976 808 5010
rect 842 4976 930 5010
rect -44 4952 68 4958
rect -44 4937 102 4952
rect -44 4919 -7 4937
rect 27 4919 102 4937
rect -44 4885 -20 4919
rect 27 4903 52 4919
rect 86 4918 102 4919
rect 14 4885 52 4903
rect -44 4884 68 4885
rect -44 4869 102 4884
rect -44 4846 -7 4869
rect 27 4850 102 4869
rect 27 4846 68 4850
rect -44 4812 -20 4846
rect 27 4835 52 4846
rect 14 4812 52 4835
rect 86 4812 102 4816
rect -44 4801 102 4812
rect -44 4773 -7 4801
rect 27 4782 102 4801
rect 27 4773 68 4782
rect -44 4739 -20 4773
rect 27 4767 52 4773
rect 14 4739 52 4767
rect 86 4739 102 4748
rect -44 4733 102 4739
rect -44 4700 -7 4733
rect 27 4714 102 4733
rect 27 4700 68 4714
rect -44 4666 -20 4700
rect 27 4699 52 4700
rect 14 4666 52 4699
rect 86 4666 102 4680
rect -44 4665 102 4666
rect -44 4631 -7 4665
rect 27 4646 102 4665
rect 27 4631 68 4646
rect -44 4627 68 4631
rect -44 4593 -20 4627
rect 14 4597 52 4627
rect 27 4593 52 4597
rect 86 4593 102 4612
rect -44 4563 -7 4593
rect 27 4578 102 4593
rect 27 4563 68 4578
rect -44 4554 68 4563
rect -44 4520 -20 4554
rect 14 4529 52 4554
rect 27 4520 52 4529
rect 86 4520 102 4544
rect -44 4495 -7 4520
rect 27 4510 102 4520
rect 27 4495 68 4510
rect -44 4481 68 4495
rect -44 4447 -20 4481
rect 14 4461 52 4481
rect 27 4447 52 4461
rect 86 4447 102 4476
rect -44 4427 -7 4447
rect 27 4442 102 4447
rect 27 4427 68 4442
rect -44 4408 68 4427
rect -44 4374 -20 4408
rect 14 4393 52 4408
rect 27 4374 52 4393
rect 86 4374 102 4408
rect -44 4359 -7 4374
rect 27 4359 68 4374
rect -44 4340 68 4359
rect -44 4335 102 4340
rect -44 4301 -20 4335
rect 14 4325 52 4335
rect 27 4301 52 4325
rect 86 4306 102 4335
rect -44 4291 -7 4301
rect 27 4291 68 4301
rect -44 4272 68 4291
rect -44 4262 102 4272
rect -44 4228 -20 4262
rect 14 4257 52 4262
rect 27 4228 52 4257
rect 86 4238 102 4262
rect -44 4223 -7 4228
rect 27 4223 68 4228
rect -44 4204 68 4223
rect -44 4189 102 4204
rect -44 4155 -20 4189
rect 27 4155 52 4189
rect 86 4170 102 4189
rect -44 4136 68 4155
rect -44 4121 102 4136
rect -44 4116 -7 4121
rect 27 4116 102 4121
rect -44 4082 -20 4116
rect 27 4087 52 4116
rect 86 4102 102 4116
rect 14 4082 52 4087
rect -44 4068 68 4082
rect -44 4053 102 4068
rect -44 4043 -7 4053
rect 27 4043 102 4053
rect -44 4009 -20 4043
rect 27 4019 52 4043
rect 86 4034 102 4043
rect 14 4009 52 4019
rect -44 4000 68 4009
rect -44 3985 102 4000
rect -44 3970 -7 3985
rect 27 3970 102 3985
rect -44 3936 -20 3970
rect 27 3951 52 3970
rect 86 3966 102 3970
rect 14 3936 52 3951
rect -44 3932 68 3936
rect -44 3917 102 3932
rect -44 3897 -7 3917
rect 27 3898 102 3917
rect 27 3897 68 3898
rect -44 3863 -20 3897
rect 27 3883 52 3897
rect 14 3863 52 3883
rect 86 3863 102 3864
rect -44 3849 102 3863
rect -44 3824 -7 3849
rect 27 3830 102 3849
rect 27 3824 68 3830
rect -44 3790 -20 3824
rect 27 3815 52 3824
rect 14 3790 52 3815
rect 86 3790 102 3796
rect -44 3781 102 3790
rect -44 3751 -7 3781
rect 27 3762 102 3781
rect 27 3751 68 3762
rect -44 3717 -20 3751
rect 27 3747 52 3751
rect 14 3717 52 3747
rect 86 3717 102 3728
rect -44 3713 102 3717
rect -44 3679 -7 3713
rect 27 3694 102 3713
rect 27 3679 68 3694
rect -44 3678 68 3679
rect -44 3644 -20 3678
rect 14 3645 52 3678
rect 27 3644 52 3645
rect 86 3644 102 3660
rect -44 3611 -7 3644
rect 27 3626 102 3644
rect 27 3611 68 3626
rect -44 3605 68 3611
rect -44 3571 -20 3605
rect 14 3577 52 3605
rect 27 3571 52 3577
rect 86 3571 102 3592
rect -44 3543 -7 3571
rect 27 3558 102 3571
rect 27 3543 68 3558
rect -44 3532 68 3543
rect -44 3498 -20 3532
rect 14 3508 52 3532
rect 27 3498 52 3508
rect 86 3498 102 3524
rect -44 3474 -7 3498
rect 27 3490 102 3498
rect 27 3474 68 3490
rect -44 3459 68 3474
rect -44 3425 -20 3459
rect 14 3439 52 3459
rect 27 3425 52 3439
rect 86 3425 102 3456
rect -44 3405 -7 3425
rect 27 3422 102 3425
rect 27 3405 68 3422
rect -44 3388 68 3405
rect -44 3386 102 3388
rect -44 3352 -20 3386
rect 14 3370 52 3386
rect 27 3352 52 3370
rect 86 3354 102 3386
rect -44 3336 -7 3352
rect 27 3336 68 3352
rect -44 3320 68 3336
rect -44 3313 102 3320
rect -44 3279 -20 3313
rect 14 3301 52 3313
rect 27 3279 52 3301
rect 86 3286 102 3313
rect -44 3267 -7 3279
rect 27 3267 68 3279
rect -44 3252 68 3267
rect -44 3240 102 3252
rect -44 3206 -20 3240
rect 14 3232 52 3240
rect 27 3206 52 3232
rect 86 3218 102 3240
rect -44 3198 -7 3206
rect 27 3198 68 3206
rect -44 3184 68 3198
rect -44 3167 102 3184
rect -44 3133 -20 3167
rect 14 3163 52 3167
rect 27 3133 52 3163
rect 86 3150 102 3167
rect -44 3129 -7 3133
rect 27 3129 68 3133
rect -44 3116 68 3129
rect -44 3094 102 3116
rect -44 3060 -20 3094
rect 27 3060 52 3094
rect 86 3082 102 3094
rect -44 3048 68 3060
rect -44 3025 102 3048
rect -44 3021 -7 3025
rect 27 3021 102 3025
rect -44 2987 -20 3021
rect 27 2991 52 3021
rect 86 3014 102 3021
rect 14 2987 52 2991
rect -44 2980 68 2987
rect -44 2956 102 2980
rect -44 2922 -7 2956
rect 27 2946 102 2956
rect 27 2922 68 2946
rect -44 2912 68 2922
rect -44 2887 102 2912
rect -44 2853 -7 2887
rect 27 2878 102 2887
rect 27 2853 68 2878
rect -44 2844 68 2853
rect -44 2818 102 2844
rect -44 2784 -7 2818
rect 27 2810 102 2818
rect 27 2784 68 2810
rect -44 2776 68 2784
rect -44 2749 102 2776
rect -44 2715 -7 2749
rect 27 2742 102 2749
rect 27 2715 68 2742
rect -44 2708 68 2715
rect -44 2704 102 2708
rect -44 2680 -3 2704
rect -44 2646 -7 2680
rect 31 2674 102 2704
rect 31 2670 68 2674
rect 27 2646 68 2670
rect -44 2640 68 2646
rect -44 2632 102 2640
rect -44 2611 -3 2632
rect -44 2577 -7 2611
rect 31 2606 102 2632
rect 31 2598 68 2606
rect 27 2577 68 2598
rect -44 2572 68 2577
rect -44 2560 102 2572
rect -44 2542 -3 2560
rect -44 2508 -7 2542
rect 31 2538 102 2560
rect 31 2526 68 2538
rect 27 2508 68 2526
rect -44 2504 68 2508
rect -44 2488 102 2504
rect -44 2473 -3 2488
rect -44 2439 -7 2473
rect 31 2470 102 2488
rect 31 2454 68 2470
rect 27 2439 68 2454
rect -44 2436 68 2439
rect -44 2416 102 2436
rect -44 2404 -3 2416
rect -44 2370 -7 2404
rect 31 2402 102 2416
rect 31 2382 68 2402
rect 27 2370 68 2382
rect -44 2368 68 2370
rect -44 2344 102 2368
rect -44 2335 -3 2344
rect -44 2301 -7 2335
rect 31 2334 102 2344
rect 31 2310 68 2334
rect 27 2301 68 2310
rect -44 2300 68 2301
rect -44 2271 102 2300
rect -44 2266 -3 2271
rect 31 2266 102 2271
rect -44 2232 -7 2266
rect 31 2237 68 2266
rect 27 2232 68 2237
rect -44 2198 102 2232
rect -44 2197 -3 2198
rect -44 2163 -7 2197
rect 31 2164 68 2198
rect 27 2163 102 2164
rect -44 2130 102 2163
rect -44 2128 68 2130
rect -44 2094 -7 2128
rect 27 2125 68 2128
rect 31 2096 68 2125
rect -44 2091 -3 2094
rect 31 2091 102 2096
rect -44 2062 102 2091
rect -44 2059 68 2062
rect -44 2025 -7 2059
rect 27 2028 68 2059
rect 27 2025 102 2028
rect -44 1994 102 2025
rect -44 1990 68 1994
rect -44 1956 -7 1990
rect 27 1960 68 1990
rect 27 1956 102 1960
rect -44 1926 102 1956
rect -44 1921 68 1926
rect -44 1887 -7 1921
rect 27 1892 68 1921
rect 27 1887 102 1892
rect -44 1858 102 1887
rect -44 1852 68 1858
rect -44 1818 -7 1852
rect 27 1824 68 1852
rect 27 1818 102 1824
rect -44 1808 102 1818
rect -10 1783 28 1808
rect -10 1774 -7 1783
rect -44 1749 -7 1774
rect 27 1774 28 1783
rect 62 1790 102 1808
rect 62 1774 68 1790
rect 27 1756 68 1774
rect 27 1749 102 1756
rect -44 1736 102 1749
rect -44 1735 28 1736
rect -10 1714 28 1735
rect -10 1701 -7 1714
rect -44 1680 -7 1701
rect 27 1702 28 1714
rect 62 1722 102 1736
rect 62 1702 68 1722
rect 27 1688 68 1702
rect 27 1680 102 1688
rect -44 1664 102 1680
rect -44 1662 28 1664
rect -10 1645 28 1662
rect -10 1628 -7 1645
rect -44 1611 -7 1628
rect 27 1630 28 1645
rect 62 1654 102 1664
rect 62 1630 68 1654
rect 27 1620 68 1630
rect 27 1611 102 1620
rect -44 1592 102 1611
rect -44 1589 28 1592
rect -10 1576 28 1589
rect -10 1555 -7 1576
rect -44 1542 -7 1555
rect 27 1558 28 1576
rect 62 1586 102 1592
rect 62 1558 68 1586
rect 27 1552 68 1558
rect 27 1542 102 1552
rect -44 1520 102 1542
rect -44 1516 28 1520
rect -10 1507 28 1516
rect -10 1482 -7 1507
rect -44 1473 -7 1482
rect 27 1486 28 1507
rect 62 1518 102 1520
rect 62 1486 68 1518
rect 27 1484 68 1486
rect 27 1473 102 1484
rect -44 1450 102 1473
rect -44 1448 68 1450
rect -44 1443 28 1448
rect -10 1438 28 1443
rect -10 1409 -7 1438
rect -44 1404 -7 1409
rect 27 1414 28 1438
rect 62 1416 68 1448
rect 62 1414 102 1416
rect 27 1404 102 1414
rect -44 1381 102 1404
rect -44 1376 68 1381
rect -44 1370 28 1376
rect -10 1369 28 1370
rect -10 1336 -7 1369
rect -44 1335 -7 1336
rect 27 1342 28 1369
rect 62 1347 68 1376
rect 62 1342 102 1347
rect 27 1335 102 1342
rect -44 1312 102 1335
rect -44 1304 68 1312
rect -44 1300 28 1304
rect -44 1297 -7 1300
rect -10 1266 -7 1297
rect 27 1270 28 1300
rect 62 1278 68 1304
rect 62 1270 102 1278
rect 27 1266 102 1270
rect -10 1263 102 1266
rect -44 1243 102 1263
rect -44 1232 68 1243
rect -44 1231 28 1232
rect -44 1224 -7 1231
rect -10 1197 -7 1224
rect 27 1198 28 1231
rect 62 1209 68 1232
rect 62 1198 102 1209
rect 27 1197 102 1198
rect -10 1190 102 1197
rect -44 1174 102 1190
rect -44 1162 68 1174
rect -44 1151 -7 1162
rect -10 1128 -7 1151
rect 27 1160 68 1162
rect 27 1128 28 1160
rect -10 1126 28 1128
rect 62 1140 68 1160
rect 62 1126 102 1140
rect -10 1117 102 1126
rect -44 1105 102 1117
rect -44 1093 68 1105
rect -44 1077 -7 1093
rect -10 1059 -7 1077
rect 27 1088 68 1093
rect 27 1059 28 1088
rect -10 1054 28 1059
rect 62 1071 68 1088
rect 62 1054 102 1071
rect -10 1043 102 1054
rect -44 1036 102 1043
rect -44 1024 68 1036
rect -44 1003 -7 1024
rect -10 990 -7 1003
rect 27 1016 68 1024
rect 27 990 28 1016
rect -10 982 28 990
rect 62 1002 68 1016
rect 62 982 102 1002
rect -10 969 102 982
rect -44 967 102 969
rect -44 955 68 967
rect -44 929 -7 955
rect -10 921 -7 929
rect 27 944 68 955
rect 27 921 28 944
rect -10 910 28 921
rect 62 933 68 944
rect 62 910 102 933
rect -10 898 102 910
rect -10 895 68 898
rect -44 886 68 895
rect -44 855 -7 886
rect -10 852 -7 855
rect 27 872 68 886
rect 27 852 28 872
rect -10 838 28 852
rect 62 864 68 872
rect 62 838 102 864
rect -10 829 102 838
rect -10 821 68 829
rect -44 817 68 821
rect -44 783 -7 817
rect 27 800 68 817
rect 27 783 28 800
rect -44 781 28 783
rect -10 766 28 781
rect 62 795 68 800
rect 62 766 102 795
rect -10 760 102 766
rect -10 748 68 760
rect -10 747 -7 748
rect -44 714 -7 747
rect 27 728 68 748
rect 27 714 28 728
rect -44 707 28 714
rect -10 694 28 707
rect 62 726 68 728
rect 62 694 102 726
rect -10 691 102 694
rect -10 679 68 691
rect -10 673 -7 679
rect -44 645 -7 673
rect 27 657 68 679
rect 27 656 102 657
rect 27 645 28 656
rect -44 633 28 645
rect -10 622 28 633
rect 62 622 102 656
rect -10 610 68 622
rect -10 599 -7 610
rect -44 576 -7 599
rect 27 588 68 610
rect 27 584 102 588
rect 27 576 28 584
rect -44 559 28 576
rect -10 550 28 559
rect 62 553 102 584
rect 62 550 68 553
rect -10 541 68 550
rect -10 525 -7 541
rect -44 507 -7 525
rect 27 519 68 541
rect 27 512 102 519
rect 27 507 28 512
rect -44 485 28 507
rect -10 478 28 485
rect 62 484 102 512
rect 62 478 68 484
rect -10 472 68 478
rect -10 451 -7 472
rect -44 438 -7 451
rect 27 450 68 472
rect 27 440 102 450
rect 27 438 28 440
rect -44 411 28 438
rect -10 406 28 411
rect 62 415 102 440
rect 62 406 68 415
rect -10 403 68 406
rect -10 377 -7 403
rect -44 369 -7 377
rect 27 381 68 403
rect 27 369 102 381
rect -44 368 102 369
rect -44 337 28 368
rect -10 334 28 337
rect 62 346 102 368
rect 62 334 68 346
rect -10 303 -7 334
rect -44 300 -7 303
rect 27 312 68 334
rect 27 300 102 312
rect -44 296 102 300
rect -44 265 28 296
rect -44 263 -7 265
rect -10 231 -7 263
rect 27 262 28 265
rect 62 277 102 296
rect 62 262 68 277
rect 27 243 68 262
rect 27 231 102 243
rect -10 229 102 231
rect -44 223 102 229
rect -44 196 28 223
rect -44 189 -7 196
rect -10 162 -7 189
rect 27 189 28 196
rect 62 208 102 223
rect 62 189 68 208
rect 27 174 68 189
rect 27 162 102 174
rect -10 155 102 162
rect -44 127 102 155
rect 154 4908 796 4924
rect 154 4900 272 4908
rect 154 4866 171 4900
rect 205 4874 272 4900
rect 306 4874 354 4908
rect 388 4874 436 4908
rect 470 4874 518 4908
rect 552 4874 601 4908
rect 635 4874 684 4908
rect 718 4874 796 4908
rect 205 4866 796 4874
rect 154 4835 796 4866
rect 154 4827 756 4835
rect 154 4793 171 4827
rect 205 4822 756 4827
rect 205 4820 278 4822
rect 312 4820 391 4822
rect 205 4793 272 4820
rect 154 4786 272 4793
rect 312 4788 351 4820
rect 306 4786 351 4788
rect 385 4788 391 4820
rect 425 4820 525 4822
rect 559 4820 756 4822
rect 425 4788 430 4820
rect 385 4786 430 4788
rect 464 4786 509 4820
rect 559 4788 588 4820
rect 543 4786 588 4788
rect 622 4798 668 4820
rect 702 4801 756 4820
rect 790 4801 796 4835
rect 622 4786 662 4798
rect 702 4786 796 4801
rect 154 4764 662 4786
rect 696 4764 796 4786
rect 154 4762 796 4764
rect 154 4758 756 4762
rect 154 4754 318 4758
rect 154 4720 171 4754
rect 205 4728 318 4754
rect 205 4720 254 4728
rect 154 4694 254 4720
rect 288 4694 318 4728
rect 523 4748 756 4758
rect 523 4729 668 4748
rect 154 4681 318 4694
rect 154 4647 171 4681
rect 205 4659 318 4681
rect 205 4647 254 4659
rect 288 4658 318 4659
rect 154 4625 254 4647
rect 154 4624 284 4625
rect 154 4608 318 4624
rect 154 4574 171 4608
rect 205 4590 318 4608
rect 205 4574 254 4590
rect 288 4583 318 4590
rect 154 4556 254 4574
rect 154 4549 284 4556
rect 154 4535 318 4549
rect 154 4501 171 4535
rect 205 4521 318 4535
rect 205 4501 254 4521
rect 288 4508 318 4521
rect 154 4487 254 4501
rect 154 4474 284 4487
rect 154 4462 318 4474
rect 154 4428 171 4462
rect 205 4452 318 4462
rect 205 4428 254 4452
rect 288 4433 318 4452
rect 154 4418 254 4428
rect 154 4399 284 4418
rect 154 4389 318 4399
rect 154 4355 171 4389
rect 205 4383 318 4389
rect 205 4355 254 4383
rect 288 4357 318 4383
rect 154 4349 254 4355
rect 154 4323 284 4349
rect 154 4315 318 4323
rect 154 4281 171 4315
rect 205 4314 318 4315
rect 205 4281 254 4314
rect 288 4281 318 4314
rect 154 4280 254 4281
rect 154 4247 284 4280
rect 154 4245 318 4247
rect 154 4241 254 4245
rect 154 4207 171 4241
rect 205 4211 254 4241
rect 288 4211 318 4245
rect 205 4207 318 4211
rect 154 4205 318 4207
rect 154 4176 284 4205
rect 154 4167 254 4176
rect 154 4133 171 4167
rect 205 4142 254 4167
rect 288 4142 318 4171
rect 205 4133 318 4142
rect 154 4129 318 4133
rect 154 4107 284 4129
rect 154 4093 254 4107
rect 154 4059 171 4093
rect 205 4073 254 4093
rect 288 4073 318 4095
rect 205 4059 318 4073
rect 154 4053 318 4059
rect 154 4038 284 4053
rect 154 4019 254 4038
rect 154 3985 171 4019
rect 205 4004 254 4019
rect 288 4004 318 4019
rect 205 3985 318 4004
rect 154 3977 318 3985
rect 154 3969 284 3977
rect 154 3945 254 3969
rect 154 3911 171 3945
rect 205 3935 254 3945
rect 288 3935 318 3943
rect 205 3911 318 3935
rect 154 3901 318 3911
rect 154 3900 284 3901
rect 154 3871 254 3900
rect 154 3837 171 3871
rect 205 3866 254 3871
rect 288 3866 318 3867
rect 205 3837 318 3866
rect 154 3831 318 3837
rect 154 3797 254 3831
rect 288 3825 318 3831
rect 154 3763 171 3797
rect 205 3791 284 3797
rect 205 3763 318 3791
rect 154 3762 318 3763
rect 154 3728 254 3762
rect 288 3728 318 3762
rect 154 3723 318 3728
rect 154 3689 171 3723
rect 205 3693 318 3723
rect 205 3689 254 3693
rect 154 3659 254 3689
rect 288 3659 318 3693
rect 154 3649 318 3659
rect 154 3615 171 3649
rect 205 3624 318 3649
rect 205 3615 254 3624
rect 154 3590 254 3615
rect 288 3590 318 3624
rect 154 3575 318 3590
rect 154 3541 171 3575
rect 205 3555 318 3575
rect 205 3541 254 3555
rect 154 3521 254 3541
rect 288 3521 318 3555
rect 154 3501 318 3521
rect 154 3467 171 3501
rect 205 3486 318 3501
rect 205 3467 254 3486
rect 154 3452 254 3467
rect 288 3452 318 3486
rect 154 3427 318 3452
rect 154 3393 171 3427
rect 205 3417 318 3427
rect 205 3393 254 3417
rect 154 3383 254 3393
rect 288 3383 318 3417
rect 154 3353 318 3383
rect 154 3319 171 3353
rect 205 3348 318 3353
rect 205 3319 254 3348
rect 154 3314 254 3319
rect 288 3314 318 3348
rect 154 3279 318 3314
rect 154 3245 171 3279
rect 205 3245 254 3279
rect 288 3245 318 3279
rect 154 3210 318 3245
rect 154 3205 254 3210
rect 154 3171 171 3205
rect 205 3176 254 3205
rect 288 3176 318 3210
rect 205 3171 318 3176
rect 154 3141 318 3171
rect 154 3131 254 3141
rect 154 3097 171 3131
rect 205 3107 254 3131
rect 288 3107 318 3141
rect 205 3097 318 3107
rect 154 3072 318 3097
rect 154 3057 254 3072
rect 154 3023 171 3057
rect 205 3038 254 3057
rect 288 3038 318 3072
rect 205 3023 318 3038
rect 154 3003 318 3023
rect 154 2969 254 3003
rect 288 2969 318 3003
rect 154 2934 318 2969
rect 154 2900 254 2934
rect 288 2900 318 2934
rect 154 2865 318 2900
rect 154 2831 254 2865
rect 288 2831 318 2865
rect 154 2796 318 2831
rect 154 2762 254 2796
rect 288 2762 318 2796
rect 154 2727 318 2762
rect 154 2702 254 2727
rect 288 2702 318 2727
rect 154 2668 164 2702
rect 198 2693 254 2702
rect 198 2668 266 2693
rect 300 2668 318 2702
rect 154 2658 318 2668
rect 154 2627 254 2658
rect 288 2627 318 2658
rect 154 2593 164 2627
rect 198 2624 254 2627
rect 198 2593 266 2624
rect 300 2593 318 2627
rect 154 2589 318 2593
rect 154 2555 254 2589
rect 288 2555 318 2589
rect 154 2551 318 2555
rect 154 2517 164 2551
rect 198 2520 266 2551
rect 198 2517 254 2520
rect 300 2517 318 2551
rect 154 2486 254 2517
rect 288 2486 318 2517
rect 154 2451 318 2486
rect 154 2417 254 2451
rect 288 2417 318 2451
rect 154 2382 318 2417
rect 154 2348 254 2382
rect 288 2348 318 2382
rect 154 2313 318 2348
rect 154 2279 254 2313
rect 288 2279 318 2313
rect 154 2270 318 2279
rect 154 2236 164 2270
rect 198 2244 266 2270
rect 198 2236 254 2244
rect 300 2236 318 2270
rect 154 2210 254 2236
rect 288 2210 318 2236
rect 154 2195 318 2210
rect 154 2161 164 2195
rect 198 2175 266 2195
rect 198 2161 254 2175
rect 300 2161 318 2195
rect 154 2141 254 2161
rect 288 2141 318 2161
rect 154 2119 318 2141
rect 154 2085 164 2119
rect 198 2106 266 2119
rect 198 2085 254 2106
rect 300 2085 318 2119
rect 154 2072 254 2085
rect 288 2072 318 2085
rect 154 2037 318 2072
rect 154 2003 254 2037
rect 288 2003 318 2037
rect 154 1968 318 2003
rect 154 1934 254 1968
rect 288 1934 318 1968
rect 154 1899 318 1934
rect 154 1865 254 1899
rect 288 1865 318 1899
rect 154 1830 318 1865
rect 154 1796 254 1830
rect 288 1796 318 1830
rect 154 1764 318 1796
rect 154 1730 167 1764
rect 201 1761 255 1764
rect 201 1730 254 1761
rect 289 1730 318 1764
rect 154 1727 254 1730
rect 288 1727 318 1730
rect 154 1692 318 1727
rect 154 1690 254 1692
rect 288 1691 318 1692
rect 154 1656 167 1690
rect 201 1658 254 1690
rect 201 1657 255 1658
rect 289 1657 318 1691
rect 201 1656 318 1657
rect 154 1623 318 1656
rect 154 1616 254 1623
rect 288 1618 318 1623
rect 154 1582 167 1616
rect 201 1589 254 1616
rect 201 1584 255 1589
rect 289 1584 318 1618
rect 201 1582 318 1584
rect 154 1554 318 1582
rect 154 1542 254 1554
rect 288 1545 318 1554
rect 154 1508 167 1542
rect 201 1520 254 1542
rect 201 1511 255 1520
rect 289 1511 318 1545
rect 201 1508 318 1511
rect 154 1485 318 1508
rect 154 1468 254 1485
rect 288 1472 318 1485
rect 154 1434 167 1468
rect 201 1451 254 1468
rect 201 1438 255 1451
rect 289 1438 318 1472
rect 201 1434 318 1438
rect 154 1416 318 1434
rect 154 1394 254 1416
rect 288 1399 318 1416
rect 154 1360 167 1394
rect 201 1382 254 1394
rect 201 1365 255 1382
rect 289 1365 318 1399
rect 201 1360 318 1365
rect 154 1347 318 1360
rect 154 1320 254 1347
rect 288 1326 318 1347
rect 154 1286 167 1320
rect 201 1313 254 1320
rect 201 1292 255 1313
rect 289 1292 318 1326
rect 201 1286 318 1292
rect 154 1278 318 1286
rect 154 1246 254 1278
rect 288 1253 318 1278
rect 154 1212 167 1246
rect 201 1244 254 1246
rect 201 1219 255 1244
rect 289 1219 318 1253
rect 201 1212 318 1219
rect 154 1209 318 1212
rect 154 1175 254 1209
rect 288 1180 318 1209
rect 154 1172 255 1175
rect 154 1138 167 1172
rect 201 1146 255 1172
rect 289 1146 318 1180
rect 201 1140 318 1146
rect 201 1138 254 1140
rect 154 1106 254 1138
rect 288 1107 318 1140
rect 154 1098 255 1106
rect 154 1064 167 1098
rect 201 1073 255 1098
rect 289 1073 318 1107
rect 201 1071 318 1073
rect 201 1064 254 1071
rect 154 1037 254 1064
rect 288 1037 318 1071
rect 154 1034 318 1037
rect 154 1025 255 1034
rect 154 991 167 1025
rect 201 1002 255 1025
rect 201 991 254 1002
rect 289 1000 318 1034
rect 154 968 254 991
rect 288 968 318 1000
rect 154 961 318 968
rect 154 952 255 961
rect 154 918 167 952
rect 201 933 255 952
rect 201 918 254 933
rect 289 927 318 961
rect 154 899 254 918
rect 288 899 318 927
rect 154 888 318 899
rect 154 879 255 888
rect 154 845 167 879
rect 201 864 255 879
rect 201 845 254 864
rect 289 854 318 888
rect 154 830 254 845
rect 288 830 318 854
rect 154 815 318 830
rect 154 806 255 815
rect 154 772 167 806
rect 201 795 255 806
rect 201 772 254 795
rect 289 781 318 815
rect 154 761 254 772
rect 288 761 318 781
rect 154 742 318 761
rect 154 733 255 742
rect 154 699 167 733
rect 201 726 255 733
rect 201 699 254 726
rect 289 708 318 742
rect 154 692 254 699
rect 288 692 318 708
rect 154 670 318 692
rect 154 660 255 670
rect 154 626 167 660
rect 201 657 255 660
rect 201 626 254 657
rect 289 636 318 670
rect 154 623 254 626
rect 288 623 318 636
rect 154 598 318 623
rect 154 588 255 598
rect 154 587 254 588
rect 154 553 167 587
rect 201 554 254 587
rect 289 564 318 598
rect 288 554 318 564
rect 201 553 318 554
rect 154 526 318 553
rect 154 519 255 526
rect 154 514 254 519
rect 154 480 167 514
rect 201 485 254 514
rect 289 492 318 526
rect 288 485 318 492
rect 201 480 318 485
rect 154 454 318 480
rect 154 450 255 454
rect 154 441 254 450
rect 154 407 167 441
rect 201 416 254 441
rect 289 420 318 454
rect 288 416 318 420
rect 201 407 318 416
rect 154 382 318 407
rect 154 381 255 382
rect 154 368 254 381
rect 154 334 167 368
rect 201 347 254 368
rect 289 348 318 382
rect 370 4702 471 4718
rect 404 4668 471 4702
rect 370 4634 471 4668
rect 404 4600 471 4634
rect 370 4566 471 4600
rect 404 4532 471 4566
rect 370 4498 471 4532
rect 404 4464 471 4498
rect 370 4430 471 4464
rect 404 4396 471 4430
rect 370 4362 471 4396
rect 404 4328 471 4362
rect 370 4294 471 4328
rect 404 4260 471 4294
rect 370 4226 471 4260
rect 404 4192 471 4226
rect 370 4158 471 4192
rect 404 4124 471 4158
rect 370 4090 471 4124
rect 404 4056 471 4090
rect 370 4022 471 4056
rect 404 3988 471 4022
rect 370 3954 471 3988
rect 404 3920 471 3954
rect 370 3886 471 3920
rect 404 3852 471 3886
rect 370 3818 471 3852
rect 404 3784 471 3818
rect 370 3725 471 3784
rect 523 4702 662 4729
rect 702 4728 756 4748
rect 790 4728 796 4762
rect 702 4714 796 4728
rect 523 4668 546 4702
rect 580 4695 662 4702
rect 696 4695 796 4714
rect 580 4689 796 4695
rect 580 4676 756 4689
rect 580 4668 668 4676
rect 523 4660 668 4668
rect 523 4658 662 4660
rect 523 4624 539 4658
rect 573 4634 662 4658
rect 702 4655 756 4676
rect 790 4655 796 4689
rect 702 4642 796 4655
rect 580 4626 662 4634
rect 696 4626 796 4642
rect 523 4600 546 4624
rect 580 4616 796 4626
rect 580 4604 756 4616
rect 580 4600 668 4604
rect 523 4591 668 4600
rect 523 4583 662 4591
rect 523 4549 539 4583
rect 573 4566 662 4583
rect 702 4582 756 4604
rect 790 4582 796 4616
rect 702 4570 796 4582
rect 580 4557 662 4566
rect 696 4557 796 4570
rect 523 4532 546 4549
rect 580 4543 796 4557
rect 580 4532 756 4543
rect 523 4522 668 4532
rect 523 4508 662 4522
rect 523 4474 539 4508
rect 573 4498 662 4508
rect 702 4509 756 4532
rect 790 4509 796 4543
rect 702 4498 796 4509
rect 580 4488 662 4498
rect 696 4488 796 4498
rect 523 4464 546 4474
rect 580 4470 796 4488
rect 580 4464 756 4470
rect 523 4459 756 4464
rect 523 4453 668 4459
rect 523 4433 662 4453
rect 523 4399 539 4433
rect 573 4430 662 4433
rect 580 4419 662 4430
rect 702 4436 756 4459
rect 790 4436 796 4470
rect 702 4425 796 4436
rect 696 4419 796 4425
rect 523 4396 546 4399
rect 580 4397 796 4419
rect 580 4396 756 4397
rect 523 4386 756 4396
rect 523 4384 668 4386
rect 523 4362 662 4384
rect 523 4357 546 4362
rect 523 4323 539 4357
rect 580 4350 662 4362
rect 702 4363 756 4386
rect 790 4363 796 4397
rect 702 4352 796 4363
rect 696 4350 796 4352
rect 580 4328 796 4350
rect 573 4324 796 4328
rect 573 4323 756 4324
rect 523 4315 756 4323
rect 523 4294 662 4315
rect 696 4313 756 4315
rect 523 4281 546 4294
rect 580 4281 662 4294
rect 702 4290 756 4313
rect 790 4290 796 4324
rect 523 4247 539 4281
rect 580 4279 668 4281
rect 702 4279 796 4290
rect 580 4260 796 4279
rect 573 4251 796 4260
rect 573 4247 756 4251
rect 523 4246 756 4247
rect 523 4226 662 4246
rect 696 4240 756 4246
rect 523 4205 546 4226
rect 580 4212 662 4226
rect 702 4217 756 4240
rect 790 4217 796 4251
rect 580 4206 668 4212
rect 702 4206 796 4217
rect 523 4171 539 4205
rect 580 4192 796 4206
rect 573 4178 796 4192
rect 573 4177 756 4178
rect 573 4171 662 4177
rect 523 4158 662 4171
rect 696 4167 756 4177
rect 523 4129 546 4158
rect 580 4143 662 4158
rect 702 4144 756 4167
rect 790 4144 796 4178
rect 580 4133 668 4143
rect 702 4133 796 4144
rect 523 4095 539 4129
rect 580 4124 796 4133
rect 573 4108 796 4124
rect 573 4095 662 4108
rect 523 4090 662 4095
rect 696 4105 796 4108
rect 696 4094 756 4105
rect 523 4056 546 4090
rect 580 4074 662 4090
rect 580 4060 668 4074
rect 702 4071 756 4094
rect 790 4071 796 4105
rect 702 4060 796 4071
rect 580 4056 796 4060
rect 523 4053 796 4056
rect 523 4019 539 4053
rect 573 4039 796 4053
rect 573 4022 662 4039
rect 523 3988 546 4019
rect 580 4005 662 4022
rect 696 4032 796 4039
rect 696 4021 756 4032
rect 580 3988 668 4005
rect 523 3987 668 3988
rect 702 3998 756 4021
rect 790 3998 796 4032
rect 702 3987 796 3998
rect 523 3977 796 3987
rect 523 3943 539 3977
rect 573 3970 796 3977
rect 573 3954 662 3970
rect 523 3920 546 3943
rect 580 3936 662 3954
rect 696 3959 796 3970
rect 696 3948 756 3959
rect 580 3920 668 3936
rect 523 3914 668 3920
rect 702 3925 756 3948
rect 790 3925 796 3959
rect 702 3914 796 3925
rect 523 3901 796 3914
rect 523 3867 539 3901
rect 573 3886 662 3901
rect 580 3867 662 3886
rect 696 3886 796 3901
rect 696 3875 756 3886
rect 523 3852 546 3867
rect 580 3852 668 3867
rect 523 3841 668 3852
rect 702 3852 756 3875
rect 790 3852 796 3886
rect 702 3841 796 3852
rect 523 3832 796 3841
rect 523 3825 662 3832
rect 523 3791 539 3825
rect 573 3818 662 3825
rect 580 3798 662 3818
rect 696 3813 796 3832
rect 696 3802 756 3813
rect 523 3784 546 3791
rect 580 3784 668 3798
rect 523 3768 668 3784
rect 702 3779 756 3802
rect 790 3779 796 3813
rect 702 3768 796 3779
rect 523 3763 796 3768
rect 523 3729 662 3763
rect 696 3740 796 3763
rect 696 3729 756 3740
rect 523 3725 668 3729
rect 370 3581 438 3725
rect 546 3695 668 3725
rect 702 3706 756 3729
rect 790 3706 796 3740
rect 702 3695 796 3706
rect 546 3694 796 3695
rect 404 3547 438 3581
rect 370 3513 438 3547
rect 404 3479 438 3513
rect 370 3467 438 3479
rect 404 3411 438 3467
rect 370 3393 438 3411
rect 404 3343 438 3393
rect 370 3319 438 3343
rect 404 3275 438 3319
rect 370 3245 438 3275
rect 404 3207 438 3245
rect 370 3173 438 3207
rect 404 3137 438 3173
rect 370 3105 438 3137
rect 404 3063 438 3105
rect 370 3037 438 3063
rect 404 2989 438 3037
rect 370 2969 438 2989
rect 404 2916 438 2969
rect 370 2901 438 2916
rect 404 2843 438 2901
rect 370 2833 438 2843
rect 404 2770 438 2833
rect 370 2765 438 2770
rect 404 2731 438 2765
rect 370 2697 438 2731
rect 404 2663 438 2697
rect 370 2460 438 2663
rect 404 2426 438 2460
rect 370 2392 438 2426
rect 404 2358 438 2392
rect 370 2324 438 2358
rect 404 2290 438 2324
rect 370 2256 438 2290
rect 404 2222 438 2256
rect 370 2188 438 2222
rect 404 2154 438 2188
rect 370 2120 438 2154
rect 404 2086 438 2120
rect 370 2052 438 2086
rect 404 2018 438 2052
rect 370 2016 438 2018
rect 404 1950 438 2016
rect 370 1942 438 1950
rect 404 1882 438 1942
rect 370 1868 438 1882
rect 404 1814 438 1868
rect 370 1794 438 1814
rect 404 1746 438 1794
rect 370 1720 438 1746
rect 404 1678 438 1720
rect 370 1646 438 1678
rect 404 1610 438 1646
rect 370 1576 438 1610
rect 404 1538 438 1576
rect 370 1498 438 1538
rect 404 1464 438 1498
rect 370 1424 438 1464
rect 404 1390 438 1424
rect 370 1350 438 1390
rect 472 3674 506 3690
rect 472 2553 506 3640
rect 472 2446 506 2519
rect 472 2374 506 2412
rect 472 1434 506 2340
rect 472 1384 506 1400
rect 546 3660 662 3694
rect 696 3667 796 3694
rect 696 3660 756 3667
rect 546 3656 756 3660
rect 546 3625 668 3656
rect 702 3633 756 3656
rect 790 3633 796 3667
rect 546 3591 662 3625
rect 702 3622 796 3633
rect 696 3593 796 3622
rect 696 3591 756 3593
rect 546 3583 756 3591
rect 546 3581 668 3583
rect 580 3556 668 3581
rect 702 3559 756 3583
rect 790 3559 796 3593
rect 580 3547 662 3556
rect 702 3549 796 3559
rect 546 3522 662 3547
rect 696 3522 796 3549
rect 546 3519 796 3522
rect 546 3513 756 3519
rect 580 3510 756 3513
rect 580 3487 668 3510
rect 580 3479 662 3487
rect 546 3453 662 3479
rect 702 3485 756 3510
rect 790 3485 796 3519
rect 702 3476 796 3485
rect 696 3453 796 3476
rect 546 3445 796 3453
rect 580 3437 756 3445
rect 580 3418 668 3437
rect 580 3411 662 3418
rect 546 3384 662 3411
rect 702 3411 756 3437
rect 790 3411 796 3445
rect 702 3403 796 3411
rect 696 3384 796 3403
rect 546 3377 796 3384
rect 580 3371 796 3377
rect 580 3364 756 3371
rect 580 3349 668 3364
rect 580 3343 662 3349
rect 546 3315 662 3343
rect 702 3337 756 3364
rect 790 3337 796 3371
rect 702 3330 796 3337
rect 696 3315 796 3330
rect 546 3309 796 3315
rect 580 3297 796 3309
rect 580 3291 756 3297
rect 580 3280 668 3291
rect 580 3275 662 3280
rect 546 3246 662 3275
rect 702 3263 756 3291
rect 790 3263 796 3297
rect 702 3257 796 3263
rect 696 3246 796 3257
rect 546 3241 796 3246
rect 580 3223 796 3241
rect 580 3218 756 3223
rect 580 3211 668 3218
rect 580 3207 662 3211
rect 546 3177 662 3207
rect 702 3189 756 3218
rect 790 3189 796 3223
rect 702 3184 796 3189
rect 696 3177 796 3184
rect 546 3173 796 3177
rect 580 3149 796 3173
rect 580 3145 756 3149
rect 580 3142 668 3145
rect 580 3139 662 3142
rect 546 3108 662 3139
rect 702 3115 756 3145
rect 790 3115 796 3149
rect 702 3111 796 3115
rect 696 3108 796 3111
rect 546 3105 796 3108
rect 580 3075 796 3105
rect 580 3073 756 3075
rect 580 3071 662 3073
rect 696 3072 756 3073
rect 546 3039 662 3071
rect 702 3041 756 3072
rect 790 3041 796 3075
rect 546 3038 668 3039
rect 702 3038 796 3041
rect 546 3037 796 3038
rect 580 3004 796 3037
rect 580 3003 662 3004
rect 546 2970 662 3003
rect 696 3001 796 3004
rect 696 2999 756 3001
rect 546 2969 668 2970
rect 580 2965 668 2969
rect 702 2967 756 2999
rect 790 2967 796 3001
rect 702 2965 796 2967
rect 580 2935 796 2965
rect 546 2901 662 2935
rect 696 2927 796 2935
rect 696 2926 756 2927
rect 580 2892 668 2901
rect 702 2893 756 2926
rect 790 2893 796 2927
rect 702 2892 796 2893
rect 580 2867 796 2892
rect 546 2866 796 2867
rect 546 2833 662 2866
rect 696 2853 796 2866
rect 580 2832 662 2833
rect 580 2819 668 2832
rect 702 2819 756 2853
rect 790 2819 796 2853
rect 580 2799 796 2819
rect 546 2797 796 2799
rect 546 2765 662 2797
rect 580 2763 662 2765
rect 696 2775 796 2797
rect 696 2763 756 2775
rect 580 2741 756 2763
rect 790 2741 796 2775
rect 580 2731 796 2741
rect 546 2728 796 2731
rect 546 2697 662 2728
rect 580 2694 662 2697
rect 696 2698 796 2728
rect 696 2694 756 2698
rect 580 2664 756 2694
rect 790 2664 796 2698
rect 580 2663 796 2664
rect 546 2659 796 2663
rect 546 2625 662 2659
rect 696 2625 796 2659
rect 546 2621 796 2625
rect 546 2590 756 2621
rect 546 2556 662 2590
rect 696 2587 756 2590
rect 790 2587 796 2621
rect 696 2556 796 2587
rect 546 2544 796 2556
rect 546 2521 756 2544
rect 546 2487 662 2521
rect 696 2510 756 2521
rect 790 2510 796 2544
rect 696 2487 796 2510
rect 546 2467 796 2487
rect 546 2460 756 2467
rect 580 2452 756 2460
rect 580 2426 662 2452
rect 546 2418 662 2426
rect 696 2433 756 2452
rect 790 2433 796 2467
rect 696 2418 796 2433
rect 546 2392 796 2418
rect 580 2390 796 2392
rect 580 2383 756 2390
rect 580 2358 662 2383
rect 546 2349 662 2358
rect 696 2356 756 2383
rect 790 2356 796 2390
rect 696 2349 796 2356
rect 546 2324 796 2349
rect 580 2314 796 2324
rect 580 2290 662 2314
rect 546 2280 662 2290
rect 696 2313 796 2314
rect 696 2280 756 2313
rect 546 2279 756 2280
rect 790 2279 796 2313
rect 546 2256 796 2279
rect 580 2245 796 2256
rect 580 2222 662 2245
rect 546 2211 662 2222
rect 696 2236 796 2245
rect 696 2211 756 2236
rect 546 2202 756 2211
rect 790 2202 796 2236
rect 546 2188 796 2202
rect 580 2176 796 2188
rect 580 2154 662 2176
rect 546 2142 662 2154
rect 696 2158 796 2176
rect 696 2142 756 2158
rect 546 2124 756 2142
rect 790 2124 796 2158
rect 546 2120 796 2124
rect 580 2107 796 2120
rect 580 2086 662 2107
rect 546 2073 662 2086
rect 696 2080 796 2107
rect 696 2073 756 2080
rect 546 2052 756 2073
rect 580 2046 756 2052
rect 790 2046 796 2080
rect 580 2038 796 2046
rect 580 2018 662 2038
rect 546 2004 662 2018
rect 696 2004 796 2038
rect 546 2002 796 2004
rect 546 1984 756 2002
rect 580 1969 756 1984
rect 580 1950 662 1969
rect 546 1935 662 1950
rect 696 1968 756 1969
rect 790 1968 796 2002
rect 696 1935 796 1968
rect 546 1924 796 1935
rect 546 1916 668 1924
rect 580 1900 668 1916
rect 580 1882 662 1900
rect 702 1890 756 1924
rect 790 1890 796 1924
rect 546 1866 662 1882
rect 696 1866 796 1890
rect 546 1851 796 1866
rect 546 1848 668 1851
rect 580 1831 668 1848
rect 702 1850 796 1851
rect 580 1814 662 1831
rect 702 1817 756 1850
rect 546 1797 662 1814
rect 696 1816 756 1817
rect 790 1816 796 1850
rect 696 1797 796 1816
rect 546 1780 796 1797
rect 580 1778 796 1780
rect 580 1762 668 1778
rect 702 1776 796 1778
rect 580 1746 662 1762
rect 546 1728 662 1746
rect 702 1744 756 1776
rect 696 1742 756 1744
rect 790 1742 796 1776
rect 696 1728 796 1742
rect 546 1712 796 1728
rect 580 1705 796 1712
rect 580 1693 668 1705
rect 702 1702 796 1705
rect 580 1678 662 1693
rect 546 1659 662 1678
rect 702 1671 756 1702
rect 696 1668 756 1671
rect 790 1668 796 1702
rect 696 1659 796 1668
rect 546 1644 796 1659
rect 580 1632 796 1644
rect 580 1624 668 1632
rect 702 1628 796 1632
rect 580 1610 662 1624
rect 546 1590 662 1610
rect 702 1598 756 1628
rect 696 1594 756 1598
rect 790 1594 796 1628
rect 696 1590 796 1594
rect 546 1576 796 1590
rect 580 1559 796 1576
rect 580 1555 668 1559
rect 580 1542 662 1555
rect 546 1521 662 1542
rect 702 1554 796 1559
rect 702 1525 756 1554
rect 696 1521 756 1525
rect 546 1520 756 1521
rect 790 1520 796 1554
rect 546 1486 796 1520
rect 546 1452 662 1486
rect 702 1480 796 1486
rect 702 1452 756 1480
rect 546 1446 756 1452
rect 790 1446 796 1480
rect 546 1417 796 1446
rect 404 1344 438 1350
rect 546 1383 662 1417
rect 696 1413 796 1417
rect 702 1406 796 1413
rect 546 1379 668 1383
rect 702 1379 756 1406
rect 546 1372 756 1379
rect 790 1372 796 1406
rect 546 1348 796 1372
rect 546 1344 662 1348
rect 404 1316 471 1344
rect 370 1292 471 1316
rect 404 1242 471 1292
rect 370 1224 471 1242
rect 404 1168 471 1224
rect 370 1156 471 1168
rect 404 1095 471 1156
rect 370 1088 471 1095
rect 404 1022 471 1088
rect 370 1020 471 1022
rect 404 986 471 1020
rect 370 983 471 986
rect 404 918 471 983
rect 370 910 471 918
rect 404 850 471 910
rect 370 837 471 850
rect 404 782 471 837
rect 370 764 471 782
rect 404 714 471 764
rect 370 680 471 714
rect 404 646 471 680
rect 370 612 471 646
rect 404 578 471 612
rect 370 544 471 578
rect 404 510 471 544
rect 370 476 471 510
rect 404 442 471 476
rect 370 408 471 442
rect 404 374 471 408
rect 370 358 471 374
rect 523 1314 662 1344
rect 696 1340 796 1348
rect 702 1332 796 1340
rect 523 1306 668 1314
rect 702 1306 756 1332
rect 523 1298 756 1306
rect 790 1298 796 1332
rect 523 1292 796 1298
rect 523 1258 546 1292
rect 580 1279 796 1292
rect 580 1258 662 1279
rect 696 1267 796 1279
rect 523 1245 662 1258
rect 702 1258 796 1267
rect 523 1233 668 1245
rect 702 1233 756 1258
rect 523 1224 756 1233
rect 790 1224 796 1258
rect 523 1190 546 1224
rect 580 1210 796 1224
rect 580 1190 662 1210
rect 696 1194 796 1210
rect 523 1176 662 1190
rect 702 1184 796 1194
rect 523 1160 668 1176
rect 702 1160 756 1184
rect 523 1156 756 1160
rect 523 1122 546 1156
rect 580 1150 756 1156
rect 790 1150 796 1184
rect 580 1141 796 1150
rect 580 1122 662 1141
rect 523 1107 662 1122
rect 696 1121 796 1141
rect 702 1110 796 1121
rect 523 1088 668 1107
rect 523 1054 546 1088
rect 580 1087 668 1088
rect 702 1087 756 1110
rect 580 1076 756 1087
rect 790 1076 796 1110
rect 580 1072 796 1076
rect 580 1054 662 1072
rect 523 1038 662 1054
rect 696 1048 796 1072
rect 523 1020 668 1038
rect 523 986 546 1020
rect 580 1014 668 1020
rect 702 1036 796 1048
rect 702 1014 756 1036
rect 580 1003 756 1014
rect 580 986 662 1003
rect 523 969 662 986
rect 696 1002 756 1003
rect 790 1002 796 1036
rect 696 975 796 1002
rect 523 952 668 969
rect 523 918 546 952
rect 580 941 668 952
rect 702 962 796 975
rect 702 941 756 962
rect 580 934 756 941
rect 580 918 662 934
rect 523 900 662 918
rect 696 928 756 934
rect 790 928 796 962
rect 696 902 796 928
rect 523 884 668 900
rect 523 850 546 884
rect 580 868 668 884
rect 702 888 796 902
rect 702 868 756 888
rect 580 865 756 868
rect 580 850 662 865
rect 523 831 662 850
rect 696 854 756 865
rect 790 854 796 888
rect 696 831 796 854
rect 523 828 796 831
rect 523 816 668 828
rect 523 782 546 816
rect 580 796 668 816
rect 702 814 796 828
rect 580 782 662 796
rect 702 794 756 814
rect 523 762 662 782
rect 696 780 756 794
rect 790 780 796 814
rect 696 762 796 780
rect 523 754 796 762
rect 523 748 668 754
rect 523 714 546 748
rect 580 727 668 748
rect 702 740 796 754
rect 580 714 662 727
rect 702 720 756 740
rect 523 693 662 714
rect 696 706 756 720
rect 790 706 796 740
rect 696 693 796 706
rect 523 680 796 693
rect 523 646 546 680
rect 580 658 668 680
rect 702 666 796 680
rect 580 646 662 658
rect 702 646 756 666
rect 523 624 662 646
rect 696 632 756 646
rect 790 632 796 666
rect 696 624 796 632
rect 523 612 796 624
rect 523 578 546 612
rect 580 606 796 612
rect 580 589 668 606
rect 702 592 796 606
rect 580 578 662 589
rect 523 555 662 578
rect 702 572 756 592
rect 696 558 756 572
rect 790 558 796 592
rect 696 555 796 558
rect 523 544 796 555
rect 523 510 546 544
rect 580 532 796 544
rect 580 520 668 532
rect 580 510 662 520
rect 523 486 662 510
rect 702 518 796 532
rect 702 498 756 518
rect 696 486 756 498
rect 523 484 756 486
rect 790 484 796 518
rect 523 476 796 484
rect 523 442 546 476
rect 580 458 796 476
rect 580 451 668 458
rect 580 442 662 451
rect 523 417 662 442
rect 702 444 796 458
rect 702 424 756 444
rect 696 417 756 424
rect 523 410 756 417
rect 790 410 796 444
rect 523 408 796 410
rect 523 374 546 408
rect 580 384 796 408
rect 580 382 668 384
rect 580 374 662 382
rect 288 347 318 348
rect 201 334 318 347
rect 154 318 318 334
rect 523 348 662 374
rect 702 369 796 384
rect 702 350 756 369
rect 696 348 756 350
rect 523 335 756 348
rect 790 335 796 369
rect 523 318 796 335
rect 154 312 796 318
rect 154 295 254 312
rect 288 310 796 312
rect 154 261 167 295
rect 201 278 254 295
rect 201 276 255 278
rect 289 276 338 310
rect 372 288 421 310
rect 455 288 504 310
rect 538 288 586 310
rect 620 288 668 310
rect 702 294 796 310
rect 386 276 421 288
rect 201 261 352 276
rect 154 254 352 261
rect 386 254 423 276
rect 457 254 494 288
rect 538 276 566 288
rect 620 276 638 288
rect 702 276 756 294
rect 528 254 566 276
rect 600 254 638 276
rect 672 260 756 276
rect 790 260 796 294
rect 672 254 796 260
rect 154 222 796 254
rect 154 188 239 222
rect 273 188 313 222
rect 347 188 387 222
rect 421 188 461 222
rect 495 188 535 222
rect 569 188 609 222
rect 643 188 683 222
rect 717 188 796 222
rect 154 154 796 188
rect -44 115 -7 127
rect -10 93 -7 115
rect 27 102 102 127
rect 848 102 930 4976
rect 27 101 92 102
rect 126 101 161 102
rect 195 101 230 102
rect 264 101 300 102
rect 334 101 370 102
rect 404 101 440 102
rect 474 101 510 102
rect 27 93 59 101
rect -10 81 59 93
rect -44 67 59 81
rect 126 68 134 101
rect 195 68 209 101
rect 264 68 284 101
rect 334 68 359 101
rect 404 68 434 101
rect 474 68 509 101
rect 544 68 580 102
rect 614 101 650 102
rect 684 101 720 102
rect 754 101 790 102
rect 824 101 930 102
rect 618 68 650 101
rect 693 68 720 101
rect 768 68 790 101
rect 93 67 134 68
rect 168 67 209 68
rect 243 67 284 68
rect 318 67 359 68
rect 393 67 434 68
rect 468 67 509 68
rect 543 67 584 68
rect 618 67 659 68
rect 693 67 734 68
rect 768 67 808 68
rect 842 67 930 101
rect -44 58 930 67
rect -44 41 -7 58
rect -10 24 -7 41
rect 27 34 930 58
rect 27 24 92 34
rect -10 7 92 24
rect -44 0 92 7
rect 126 0 161 34
rect 195 0 230 34
rect 264 0 300 34
rect 334 0 370 34
rect 404 0 440 34
rect 474 0 510 34
rect 544 0 580 34
rect 614 0 650 34
rect 684 0 720 34
rect 754 0 790 34
rect 824 0 930 34
rect -44 -34 930 0
rect 848 -36 930 -34
<< viali >>
rect -20 12111 -7 12129
rect -7 12111 14 12129
rect -20 12095 14 12111
rect 52 12095 86 12129
rect -20 12043 -7 12055
rect -7 12043 14 12055
rect -20 12021 14 12043
rect 52 12021 86 12055
rect 163 12010 197 12044
rect 246 12010 280 12044
rect 329 12010 363 12044
rect 412 12010 446 12044
rect 496 12010 530 12044
rect 580 12010 614 12044
rect 664 12010 698 12044
rect -20 11975 -7 11981
rect -7 11975 14 11981
rect -20 11947 14 11975
rect 52 11947 86 11981
rect -20 11873 14 11907
rect 52 11873 86 11907
rect -20 11805 14 11833
rect -20 11799 -7 11805
rect -7 11799 14 11805
rect 52 11799 86 11833
rect -20 11737 14 11759
rect -20 11725 -7 11737
rect -7 11725 14 11737
rect 52 11725 86 11759
rect -20 11669 14 11685
rect -20 11651 -7 11669
rect -7 11651 14 11669
rect 52 11651 86 11685
rect -20 11601 14 11611
rect -20 11577 -7 11601
rect -7 11577 14 11601
rect 52 11577 86 11611
rect -20 11533 14 11537
rect -20 11503 -7 11533
rect -7 11503 14 11533
rect 52 11503 86 11537
rect -20 11431 -7 11463
rect -7 11431 14 11463
rect -20 11429 14 11431
rect 52 11429 86 11463
rect -20 11363 -7 11389
rect -7 11363 14 11389
rect -20 11355 14 11363
rect 52 11355 86 11389
rect -20 11295 -7 11315
rect -7 11295 14 11315
rect -20 11281 14 11295
rect 52 11281 86 11315
rect -20 11227 -7 11241
rect -7 11227 14 11241
rect -20 11207 14 11227
rect 52 11207 86 11241
rect -20 11159 -7 11167
rect -7 11159 14 11167
rect -20 11133 14 11159
rect 52 11133 86 11167
rect -20 11091 -7 11093
rect -7 11091 14 11093
rect -20 11059 14 11091
rect 52 11059 86 11093
rect -20 10989 14 11019
rect -20 10985 -7 10989
rect -7 10985 14 10989
rect 52 10985 86 11019
rect -20 10921 14 10945
rect -20 10911 -7 10921
rect -7 10911 14 10921
rect 52 10911 86 10945
rect -20 10853 14 10871
rect -20 10837 -7 10853
rect -7 10837 14 10853
rect 52 10837 86 10871
rect -20 10785 14 10797
rect -20 10763 -7 10785
rect -7 10763 14 10785
rect 52 10763 86 10797
rect -20 10717 14 10723
rect -20 10689 -7 10717
rect -7 10689 14 10717
rect 52 10689 86 10723
rect -20 10615 -7 10649
rect -7 10615 14 10649
rect 52 10615 86 10649
rect -20 10547 -7 10575
rect -7 10547 14 10575
rect -20 10541 14 10547
rect 52 10541 86 10575
rect -20 10479 -7 10502
rect -7 10479 14 10502
rect -20 10468 14 10479
rect 52 10468 86 10502
rect 230 11925 264 11959
rect 302 11925 336 11959
rect 374 11925 408 11959
rect 446 11925 480 11959
rect 518 11925 552 11959
rect 590 11925 624 11959
rect 158 11853 192 11887
rect 158 11777 192 11811
rect 158 11701 192 11735
rect 158 11625 192 11659
rect 158 11549 192 11583
rect 158 11473 192 11507
rect 158 11397 192 11431
rect 158 11321 192 11355
rect 158 11245 192 11279
rect 158 11169 192 11203
rect 158 11093 192 11127
rect 158 11017 192 11051
rect 158 10941 192 10975
rect 158 10865 192 10899
rect 158 10789 192 10823
rect 158 10713 192 10747
rect 158 10638 192 10672
rect 158 10563 192 10597
rect 158 10488 192 10522
rect 662 11853 696 11887
rect 662 11781 696 11815
rect 662 11709 696 11743
rect 662 11637 696 11671
rect 662 11565 696 11599
rect 662 11493 696 11527
rect 662 11421 696 11455
rect 662 11349 696 11383
rect 662 11277 696 11311
rect 662 11205 696 11239
rect 662 11133 696 11167
rect 662 11061 696 11095
rect 662 10989 696 11023
rect 662 10917 696 10951
rect 662 10845 696 10879
rect 662 10773 696 10807
rect 662 10701 696 10735
rect 662 10629 696 10663
rect 662 10557 696 10591
rect 662 10485 696 10519
rect -20 10411 -7 10429
rect -7 10411 14 10429
rect -20 10395 14 10411
rect 52 10395 86 10429
rect -20 10343 -7 10356
rect -7 10343 14 10356
rect -20 10322 14 10343
rect 52 10322 86 10356
rect -20 10275 -7 10283
rect -7 10275 14 10283
rect -20 10249 14 10275
rect 52 10249 86 10283
rect -20 10207 -7 10210
rect -7 10207 14 10210
rect -20 10176 14 10207
rect 52 10176 86 10210
rect -20 10105 14 10137
rect -20 10103 -7 10105
rect -7 10103 14 10105
rect 52 10103 86 10137
rect -20 10037 14 10064
rect -20 10030 -7 10037
rect -7 10030 14 10037
rect 52 10030 86 10064
rect -20 9969 14 9991
rect -20 9957 -7 9969
rect -7 9957 14 9969
rect 52 9957 86 9991
rect -20 9901 14 9918
rect -20 9884 -7 9901
rect -7 9884 14 9901
rect 52 9884 86 9918
rect 158 10405 192 10439
rect 278 10405 312 10439
rect 158 10326 192 10360
rect 278 10326 312 10360
rect 158 10247 192 10281
rect 278 10247 312 10281
rect 158 10168 192 10202
rect 278 10168 312 10202
rect 158 10089 192 10123
rect 278 10089 312 10123
rect 158 10009 192 10043
rect 278 10009 312 10043
rect 158 9929 192 9963
rect 278 9929 312 9963
rect 158 9849 192 9883
rect 278 9849 312 9883
rect 662 10413 696 10447
rect 662 10341 696 10375
rect 662 10269 696 10303
rect 662 10197 696 10231
rect 662 10125 696 10159
rect 662 10053 696 10087
rect 662 9981 696 10015
rect 662 9909 696 9943
rect -20 9833 14 9845
rect -20 9811 -7 9833
rect -7 9811 14 9833
rect 52 9811 86 9845
rect -20 9765 14 9772
rect -20 9738 -7 9765
rect -7 9738 14 9765
rect 52 9738 86 9772
rect -20 9697 14 9699
rect -20 9665 -7 9697
rect -7 9665 14 9697
rect 52 9665 86 9699
rect -20 9595 -7 9626
rect -7 9595 14 9626
rect -20 9592 14 9595
rect 52 9592 86 9626
rect -20 9527 -7 9553
rect -7 9527 14 9553
rect -20 9519 14 9527
rect 52 9519 86 9553
rect -20 9459 -7 9480
rect -7 9459 14 9480
rect -20 9446 14 9459
rect 52 9446 86 9480
rect 662 9837 696 9871
rect 662 9765 696 9799
rect 662 9693 696 9727
rect 662 9621 696 9655
rect 662 9549 696 9583
rect 662 9477 696 9511
rect 662 9405 696 9439
rect 662 9333 696 9367
rect 662 9260 696 9294
rect 662 9187 696 9221
rect -20 9153 14 9163
rect -20 9129 -7 9153
rect -7 9129 14 9153
rect 52 9129 86 9163
rect -20 9085 14 9088
rect -20 9054 -7 9085
rect -7 9054 14 9085
rect 52 9054 86 9088
rect -20 8983 -7 9013
rect -7 8983 14 9013
rect -20 8979 14 8983
rect 52 8979 86 9013
rect -20 8915 -7 8938
rect -7 8915 14 8938
rect -20 8904 14 8915
rect 52 8904 86 8938
rect -20 8847 -7 8863
rect -7 8847 14 8863
rect -20 8829 14 8847
rect 52 8829 86 8863
rect -20 8779 -7 8788
rect -7 8779 14 8788
rect -20 8754 14 8779
rect 52 8754 86 8788
rect -20 8711 -7 8713
rect -7 8711 14 8713
rect -20 8679 14 8711
rect 52 8679 86 8713
rect -20 8609 14 8638
rect -20 8604 -7 8609
rect -7 8604 14 8609
rect 52 8604 86 8638
rect 662 9114 696 9148
rect 662 9041 696 9075
rect 662 8968 696 9002
rect 662 8895 696 8929
rect 662 8822 696 8856
rect 662 8749 696 8783
rect 662 8676 696 8710
rect -20 8541 14 8563
rect -20 8529 -7 8541
rect -7 8529 14 8541
rect 52 8529 86 8563
rect -20 8473 14 8488
rect -20 8454 -7 8473
rect -7 8454 14 8473
rect 52 8454 86 8488
rect -20 8405 14 8413
rect -20 8379 -7 8405
rect -7 8379 14 8405
rect 52 8379 86 8413
rect -20 8337 14 8338
rect -20 8304 -7 8337
rect -7 8304 14 8337
rect 52 8304 86 8338
rect -20 8235 -7 8263
rect -7 8235 14 8263
rect -20 8229 14 8235
rect 52 8229 86 8263
rect -20 8167 -7 8188
rect -7 8167 14 8188
rect -20 8154 14 8167
rect 52 8154 86 8188
rect -20 8099 -7 8113
rect -7 8099 14 8113
rect -20 8079 14 8099
rect 52 8079 86 8113
rect -20 8031 -7 8038
rect -7 8031 14 8038
rect -20 8004 14 8031
rect 52 8004 86 8038
rect 158 8587 192 8621
rect 278 8587 312 8621
rect 158 8508 192 8542
rect 278 8508 312 8542
rect 158 8429 192 8463
rect 278 8429 312 8463
rect 158 8350 192 8384
rect 278 8350 312 8384
rect 158 8271 192 8305
rect 278 8271 312 8305
rect 158 8191 192 8225
rect 278 8191 312 8225
rect 158 8111 192 8145
rect 278 8111 312 8145
rect 158 8031 192 8065
rect 278 8031 312 8065
rect 662 8603 696 8637
rect 662 8530 696 8564
rect 662 8457 696 8491
rect 662 8384 696 8418
rect 662 8311 696 8345
rect 662 8238 696 8272
rect 662 8165 696 8199
rect 662 8092 696 8126
rect -20 7929 14 7963
rect 52 7929 86 7963
rect -20 7861 14 7889
rect -20 7855 -7 7861
rect -7 7855 14 7861
rect 52 7855 86 7889
rect -20 7793 14 7815
rect -20 7781 -7 7793
rect -7 7781 14 7793
rect 52 7781 86 7815
rect -20 7725 14 7741
rect -20 7707 -7 7725
rect -7 7707 14 7725
rect 52 7707 86 7741
rect -20 7657 14 7667
rect -20 7633 -7 7657
rect -7 7633 14 7657
rect 52 7633 86 7667
rect -20 7589 14 7593
rect -20 7559 -7 7589
rect -7 7559 14 7589
rect 52 7559 86 7593
rect 662 8019 696 8053
rect 662 7946 696 7980
rect 662 7873 696 7907
rect 662 7800 696 7834
rect 662 7727 696 7761
rect 662 7654 696 7688
rect 662 7581 696 7615
rect 662 7508 696 7542
rect 662 7435 696 7469
rect 662 7362 696 7396
rect 662 7289 696 7323
rect -20 7249 14 7268
rect -20 7234 -7 7249
rect -7 7234 14 7249
rect 52 7234 86 7268
rect -20 7181 14 7194
rect -20 7160 -7 7181
rect -7 7160 14 7181
rect 52 7160 86 7194
rect -20 7113 14 7120
rect -20 7086 -7 7113
rect -7 7086 14 7113
rect 52 7086 86 7120
rect -20 7045 14 7046
rect -20 7012 -7 7045
rect -7 7012 14 7045
rect 52 7012 86 7046
rect -20 6943 -7 6972
rect -7 6943 14 6972
rect -20 6938 14 6943
rect 52 6938 86 6972
rect -20 6875 -7 6898
rect -7 6875 14 6898
rect -20 6864 14 6875
rect 52 6864 86 6898
rect -20 6807 -7 6824
rect -7 6807 14 6824
rect -20 6790 14 6807
rect 52 6790 86 6824
rect -20 6739 -7 6750
rect -7 6739 14 6750
rect -20 6716 14 6739
rect 52 6716 86 6750
rect -20 6671 -7 6676
rect -7 6671 14 6676
rect -20 6642 14 6671
rect 52 6642 86 6676
rect -20 6569 14 6602
rect -20 6568 -7 6569
rect -7 6568 14 6569
rect 52 6568 86 6602
rect -20 6501 14 6528
rect -20 6494 -7 6501
rect -7 6494 14 6501
rect 52 6494 86 6528
rect -20 6433 14 6454
rect -20 6420 -7 6433
rect -7 6420 14 6433
rect 52 6420 86 6454
rect -20 6365 14 6380
rect -20 6346 -7 6365
rect -7 6346 14 6365
rect 52 6346 86 6380
rect -20 6297 14 6306
rect -20 6272 -7 6297
rect -7 6272 14 6297
rect 52 6272 86 6306
rect -20 6229 14 6233
rect -20 6199 -7 6229
rect -7 6199 14 6229
rect 52 6199 86 6233
rect -20 6127 -7 6160
rect -7 6127 14 6160
rect -20 6126 14 6127
rect 52 6126 86 6160
rect -20 6059 -7 6087
rect -7 6059 14 6087
rect -20 6053 14 6059
rect 52 6053 86 6087
rect -20 5991 -7 6014
rect -7 5991 14 6014
rect -20 5980 14 5991
rect 52 5980 86 6014
rect -20 5923 -7 5941
rect -7 5923 14 5941
rect -20 5907 14 5923
rect 52 5907 86 5941
rect -20 5855 -7 5868
rect -7 5855 14 5868
rect -20 5834 14 5855
rect 52 5834 86 5868
rect -20 5787 -7 5795
rect -7 5787 14 5795
rect -20 5761 14 5787
rect 52 5761 86 5795
rect -20 5719 -7 5722
rect -7 5719 14 5722
rect -20 5688 14 5719
rect 52 5688 86 5722
rect -20 5617 14 5649
rect -20 5615 -7 5617
rect -7 5615 14 5617
rect 52 5615 86 5649
rect -20 5549 14 5576
rect -20 5542 -7 5549
rect -7 5542 14 5549
rect 52 5542 86 5576
rect -20 5481 14 5503
rect -20 5469 -7 5481
rect -7 5469 14 5481
rect 52 5469 86 5503
rect -20 5413 14 5430
rect -20 5396 -7 5413
rect -7 5396 14 5413
rect 52 5396 86 5430
rect -20 5345 14 5357
rect -20 5323 -7 5345
rect -7 5323 14 5345
rect 52 5323 86 5357
rect -20 5277 14 5284
rect -20 5250 -7 5277
rect -7 5250 14 5277
rect 52 5250 86 5284
rect -20 5209 14 5211
rect -20 5177 -7 5209
rect -7 5177 14 5209
rect 52 5177 86 5211
rect -20 5107 -7 5138
rect -7 5107 14 5138
rect -20 5104 14 5107
rect 52 5104 86 5138
rect 171 7239 205 7273
rect 171 7165 205 7199
rect 171 7091 205 7125
rect 171 7018 205 7052
rect 171 6945 205 6979
rect 171 6872 205 6906
rect 171 6799 205 6833
rect 171 6726 205 6760
rect 171 6653 205 6687
rect 171 6580 205 6614
rect 171 6507 205 6541
rect 171 6434 205 6468
rect 171 6361 205 6395
rect 171 6288 205 6322
rect 171 6215 205 6249
rect 171 6142 205 6176
rect 171 6069 205 6103
rect 171 5996 205 6030
rect 171 5923 205 5957
rect 171 5850 205 5884
rect 171 5777 205 5811
rect 171 5704 205 5738
rect 171 5631 205 5665
rect 171 5558 205 5592
rect 171 5485 205 5519
rect 171 5412 205 5446
rect 171 5339 205 5373
rect 171 5266 205 5300
rect 171 5193 205 5227
rect 662 7216 696 7250
rect 662 7143 696 7177
rect 662 7070 696 7104
rect 662 6997 696 7031
rect 662 6924 696 6958
rect 662 6851 696 6885
rect 662 6778 696 6812
rect 662 6705 696 6739
rect 662 6632 696 6666
rect 662 6559 696 6593
rect 662 6486 696 6520
rect 662 6413 696 6447
rect 662 6340 696 6374
rect 662 6267 696 6301
rect 662 6194 696 6228
rect 662 6121 696 6155
rect 662 6048 696 6082
rect 662 5975 696 6009
rect 662 5902 696 5936
rect 662 5829 696 5863
rect 662 5756 696 5790
rect 662 5683 696 5717
rect 662 5610 696 5644
rect 662 5537 696 5571
rect 662 5464 696 5498
rect 662 5391 696 5425
rect 662 5318 696 5352
rect 662 5245 696 5279
rect 297 5173 331 5207
rect 370 5173 404 5207
rect 443 5173 477 5207
rect 516 5173 550 5207
rect 589 5173 623 5207
rect 736 11938 770 11972
rect 736 11866 770 11900
rect 736 11794 770 11828
rect 736 11722 770 11756
rect 736 11650 770 11684
rect 736 11578 770 11612
rect 736 11506 770 11540
rect 736 11434 770 11468
rect 736 11362 770 11396
rect 736 11290 770 11324
rect 736 11218 770 11252
rect 736 11146 770 11180
rect 736 11074 770 11108
rect 736 11002 770 11036
rect 736 10930 770 10964
rect 736 10858 770 10892
rect 736 10786 770 10820
rect 736 10714 770 10748
rect 736 10642 770 10676
rect 736 10570 770 10604
rect 736 10498 770 10532
rect 736 10426 770 10460
rect 736 10354 770 10388
rect 736 10282 770 10316
rect 736 10210 770 10244
rect 736 10138 770 10172
rect 736 10066 770 10100
rect 736 9994 770 10028
rect 736 9922 770 9956
rect 736 9850 770 9884
rect 736 9778 770 9812
rect 736 9706 770 9740
rect 736 9634 770 9668
rect 736 9562 770 9596
rect 736 9490 770 9524
rect 736 9418 770 9452
rect 736 9346 770 9380
rect 736 9274 770 9308
rect 736 9202 770 9236
rect 736 9130 770 9164
rect 736 9058 770 9092
rect 736 8986 770 9020
rect 736 8914 770 8948
rect 736 8842 770 8876
rect 736 8770 770 8804
rect 736 8698 770 8732
rect 736 8626 770 8660
rect 736 8554 770 8588
rect 736 8482 770 8516
rect 736 8410 770 8444
rect 736 8338 770 8372
rect 736 8266 770 8300
rect 736 8194 770 8228
rect 736 8122 770 8156
rect 736 8050 770 8084
rect 736 7978 770 8012
rect 736 7906 770 7940
rect 736 7834 770 7868
rect 736 7762 770 7796
rect 736 7690 770 7724
rect 736 7618 770 7652
rect 736 7546 770 7580
rect 736 7474 770 7508
rect 736 7402 770 7436
rect 736 7330 770 7364
rect 736 7258 770 7292
rect 736 7186 770 7220
rect 736 7114 770 7148
rect 736 7042 770 7076
rect 736 6970 770 7004
rect 736 6898 770 6932
rect 736 6826 770 6860
rect 736 6754 770 6788
rect 736 6682 770 6716
rect 736 6610 770 6644
rect 736 6538 770 6572
rect 736 6466 770 6500
rect 736 6394 770 6428
rect 736 6322 770 6356
rect 736 6250 770 6284
rect 736 6178 770 6212
rect 736 6106 770 6140
rect 736 6034 770 6068
rect 736 5962 770 5996
rect 736 5890 770 5924
rect 736 5818 770 5852
rect 736 5746 770 5780
rect 736 5674 770 5708
rect 736 5602 770 5636
rect 736 5530 770 5564
rect 736 5458 770 5492
rect 736 5386 770 5420
rect 736 5314 770 5348
rect 736 5241 770 5275
rect 171 5120 205 5154
rect 736 5168 770 5202
rect 297 5096 331 5130
rect 371 5096 405 5130
rect 444 5096 478 5130
rect 517 5096 551 5130
rect 590 5096 624 5130
rect 663 5096 697 5130
rect -20 5039 -7 5065
rect -7 5039 14 5065
rect -20 5031 14 5039
rect 52 5031 86 5065
rect -20 4971 -7 4992
rect -7 4971 14 4992
rect 52 4986 86 4992
rect -20 4958 14 4971
rect 52 4958 68 4986
rect 68 4958 86 4986
rect 129 4976 163 5010
rect 205 4976 239 5010
rect 281 4976 315 5010
rect 357 4976 391 5010
rect 433 4976 467 5010
rect 508 4976 542 5010
rect 583 4976 617 5010
rect 658 4976 692 5010
rect 733 4976 767 5010
rect 808 4976 842 5010
rect -20 4903 -7 4919
rect -7 4903 14 4919
rect 52 4918 86 4919
rect -20 4885 14 4903
rect 52 4885 68 4918
rect 68 4885 86 4918
rect -20 4835 -7 4846
rect -7 4835 14 4846
rect -20 4812 14 4835
rect 52 4816 68 4846
rect 68 4816 86 4846
rect 52 4812 86 4816
rect -20 4767 -7 4773
rect -7 4767 14 4773
rect -20 4739 14 4767
rect 52 4748 68 4773
rect 68 4748 86 4773
rect 52 4739 86 4748
rect -20 4699 -7 4700
rect -7 4699 14 4700
rect -20 4666 14 4699
rect 52 4680 68 4700
rect 68 4680 86 4700
rect 52 4666 86 4680
rect -20 4597 14 4627
rect 52 4612 68 4627
rect 68 4612 86 4627
rect -20 4593 -7 4597
rect -7 4593 14 4597
rect 52 4593 86 4612
rect -20 4529 14 4554
rect 52 4544 68 4554
rect 68 4544 86 4554
rect -20 4520 -7 4529
rect -7 4520 14 4529
rect 52 4520 86 4544
rect -20 4461 14 4481
rect 52 4476 68 4481
rect 68 4476 86 4481
rect -20 4447 -7 4461
rect -7 4447 14 4461
rect 52 4447 86 4476
rect -20 4393 14 4408
rect -20 4374 -7 4393
rect -7 4374 14 4393
rect 52 4374 86 4408
rect -20 4325 14 4335
rect -20 4301 -7 4325
rect -7 4301 14 4325
rect 52 4306 86 4335
rect 52 4301 68 4306
rect 68 4301 86 4306
rect -20 4257 14 4262
rect -20 4228 -7 4257
rect -7 4228 14 4257
rect 52 4238 86 4262
rect 52 4228 68 4238
rect 68 4228 86 4238
rect -20 4155 -7 4189
rect -7 4155 14 4189
rect 52 4170 86 4189
rect 52 4155 68 4170
rect 68 4155 86 4170
rect -20 4087 -7 4116
rect -7 4087 14 4116
rect 52 4102 86 4116
rect -20 4082 14 4087
rect 52 4082 68 4102
rect 68 4082 86 4102
rect -20 4019 -7 4043
rect -7 4019 14 4043
rect 52 4034 86 4043
rect -20 4009 14 4019
rect 52 4009 68 4034
rect 68 4009 86 4034
rect -20 3951 -7 3970
rect -7 3951 14 3970
rect 52 3966 86 3970
rect -20 3936 14 3951
rect 52 3936 68 3966
rect 68 3936 86 3966
rect -20 3883 -7 3897
rect -7 3883 14 3897
rect -20 3863 14 3883
rect 52 3864 68 3897
rect 68 3864 86 3897
rect 52 3863 86 3864
rect -20 3815 -7 3824
rect -7 3815 14 3824
rect -20 3790 14 3815
rect 52 3796 68 3824
rect 68 3796 86 3824
rect 52 3790 86 3796
rect -20 3747 -7 3751
rect -7 3747 14 3751
rect -20 3717 14 3747
rect 52 3728 68 3751
rect 68 3728 86 3751
rect 52 3717 86 3728
rect -20 3645 14 3678
rect 52 3660 68 3678
rect 68 3660 86 3678
rect -20 3644 -7 3645
rect -7 3644 14 3645
rect 52 3644 86 3660
rect -20 3577 14 3605
rect 52 3592 68 3605
rect 68 3592 86 3605
rect -20 3571 -7 3577
rect -7 3571 14 3577
rect 52 3571 86 3592
rect -20 3508 14 3532
rect 52 3524 68 3532
rect 68 3524 86 3532
rect -20 3498 -7 3508
rect -7 3498 14 3508
rect 52 3498 86 3524
rect -20 3439 14 3459
rect 52 3456 68 3459
rect 68 3456 86 3459
rect -20 3425 -7 3439
rect -7 3425 14 3439
rect 52 3425 86 3456
rect -20 3370 14 3386
rect -20 3352 -7 3370
rect -7 3352 14 3370
rect 52 3354 86 3386
rect 52 3352 68 3354
rect 68 3352 86 3354
rect -20 3301 14 3313
rect -20 3279 -7 3301
rect -7 3279 14 3301
rect 52 3286 86 3313
rect 52 3279 68 3286
rect 68 3279 86 3286
rect -20 3232 14 3240
rect -20 3206 -7 3232
rect -7 3206 14 3232
rect 52 3218 86 3240
rect 52 3206 68 3218
rect 68 3206 86 3218
rect -20 3163 14 3167
rect -20 3133 -7 3163
rect -7 3133 14 3163
rect 52 3150 86 3167
rect 52 3133 68 3150
rect 68 3133 86 3150
rect -20 3060 -7 3094
rect -7 3060 14 3094
rect 52 3082 86 3094
rect 52 3060 68 3082
rect 68 3060 86 3082
rect -20 2991 -7 3021
rect -7 2991 14 3021
rect 52 3014 86 3021
rect -20 2987 14 2991
rect 52 2987 68 3014
rect 68 2987 86 3014
rect -3 2680 31 2704
rect -3 2670 27 2680
rect 27 2670 31 2680
rect -3 2611 31 2632
rect -3 2598 27 2611
rect 27 2598 31 2611
rect -3 2542 31 2560
rect -3 2526 27 2542
rect 27 2526 31 2542
rect -3 2473 31 2488
rect -3 2454 27 2473
rect 27 2454 31 2473
rect -3 2404 31 2416
rect -3 2382 27 2404
rect 27 2382 31 2404
rect -3 2335 31 2344
rect -3 2310 27 2335
rect 27 2310 31 2335
rect -3 2266 31 2271
rect -3 2237 27 2266
rect 27 2237 31 2266
rect -3 2197 31 2198
rect -3 2164 27 2197
rect 27 2164 31 2197
rect -3 2094 27 2125
rect 27 2094 31 2125
rect -3 2091 31 2094
rect -44 1774 -10 1808
rect 28 1774 62 1808
rect -44 1701 -10 1735
rect 28 1702 62 1736
rect -44 1628 -10 1662
rect 28 1630 62 1664
rect -44 1555 -10 1589
rect 28 1558 62 1592
rect -44 1482 -10 1516
rect 28 1486 62 1520
rect -44 1409 -10 1443
rect 28 1414 62 1448
rect -44 1336 -10 1370
rect 28 1342 62 1376
rect -44 1263 -10 1297
rect 28 1270 62 1304
rect -44 1190 -10 1224
rect 28 1198 62 1232
rect -44 1117 -10 1151
rect 28 1126 62 1160
rect -44 1043 -10 1077
rect 28 1054 62 1088
rect -44 969 -10 1003
rect 28 982 62 1016
rect -44 895 -10 929
rect 28 910 62 944
rect -44 821 -10 855
rect 28 838 62 872
rect -44 747 -10 781
rect 28 766 62 800
rect -44 673 -10 707
rect 28 694 62 728
rect -44 599 -10 633
rect 28 622 62 656
rect -44 525 -10 559
rect 28 550 62 584
rect -44 451 -10 485
rect 28 478 62 512
rect -44 377 -10 411
rect 28 406 62 440
rect -44 303 -10 337
rect 28 334 62 368
rect -44 229 -10 263
rect 28 262 62 296
rect -44 155 -10 189
rect 28 189 62 223
rect 171 4866 205 4900
rect 272 4874 306 4908
rect 354 4874 388 4908
rect 436 4874 470 4908
rect 518 4874 552 4908
rect 601 4874 635 4908
rect 684 4874 718 4908
rect 171 4793 205 4827
rect 272 4788 278 4820
rect 278 4788 306 4820
rect 272 4786 306 4788
rect 351 4786 385 4820
rect 430 4786 464 4820
rect 509 4788 525 4820
rect 525 4788 543 4820
rect 509 4786 543 4788
rect 588 4786 622 4820
rect 668 4798 702 4820
rect 756 4801 790 4835
rect 668 4786 696 4798
rect 696 4786 702 4798
rect 171 4720 205 4754
rect 668 4729 702 4748
rect 171 4647 205 4681
rect 284 4625 288 4658
rect 288 4625 318 4658
rect 284 4624 318 4625
rect 171 4574 205 4608
rect 284 4556 288 4583
rect 288 4556 318 4583
rect 284 4549 318 4556
rect 171 4501 205 4535
rect 284 4487 288 4508
rect 288 4487 318 4508
rect 284 4474 318 4487
rect 171 4428 205 4462
rect 284 4418 288 4433
rect 288 4418 318 4433
rect 284 4399 318 4418
rect 171 4355 205 4389
rect 284 4349 288 4357
rect 288 4349 318 4357
rect 284 4323 318 4349
rect 171 4281 205 4315
rect 284 4280 288 4281
rect 288 4280 318 4281
rect 284 4247 318 4280
rect 171 4207 205 4241
rect 284 4176 318 4205
rect 284 4171 288 4176
rect 288 4171 318 4176
rect 171 4133 205 4167
rect 284 4107 318 4129
rect 284 4095 288 4107
rect 288 4095 318 4107
rect 171 4059 205 4093
rect 284 4038 318 4053
rect 284 4019 288 4038
rect 288 4019 318 4038
rect 171 3985 205 4019
rect 284 3969 318 3977
rect 171 3911 205 3945
rect 284 3943 288 3969
rect 288 3943 318 3969
rect 284 3900 318 3901
rect 171 3837 205 3871
rect 284 3867 288 3900
rect 288 3867 318 3900
rect 284 3797 288 3825
rect 288 3797 318 3825
rect 171 3763 205 3797
rect 284 3791 318 3797
rect 171 3689 205 3723
rect 171 3615 205 3649
rect 171 3541 205 3575
rect 171 3467 205 3501
rect 171 3393 205 3427
rect 171 3319 205 3353
rect 171 3245 205 3279
rect 171 3171 205 3205
rect 171 3097 205 3131
rect 171 3023 205 3057
rect 164 2668 198 2702
rect 266 2693 288 2702
rect 288 2693 300 2702
rect 266 2668 300 2693
rect 164 2593 198 2627
rect 266 2624 288 2627
rect 288 2624 300 2627
rect 266 2593 300 2624
rect 164 2517 198 2551
rect 266 2520 300 2551
rect 266 2517 288 2520
rect 288 2517 300 2520
rect 164 2236 198 2270
rect 266 2244 300 2270
rect 266 2236 288 2244
rect 288 2236 300 2244
rect 164 2161 198 2195
rect 266 2175 300 2195
rect 266 2161 288 2175
rect 288 2161 300 2175
rect 164 2085 198 2119
rect 266 2106 300 2119
rect 266 2085 288 2106
rect 288 2085 300 2106
rect 167 1730 201 1764
rect 255 1761 289 1764
rect 255 1730 288 1761
rect 288 1730 289 1761
rect 167 1656 201 1690
rect 255 1658 288 1691
rect 288 1658 289 1691
rect 255 1657 289 1658
rect 167 1582 201 1616
rect 255 1589 288 1618
rect 288 1589 289 1618
rect 255 1584 289 1589
rect 167 1508 201 1542
rect 255 1520 288 1545
rect 288 1520 289 1545
rect 255 1511 289 1520
rect 167 1434 201 1468
rect 255 1451 288 1472
rect 288 1451 289 1472
rect 255 1438 289 1451
rect 167 1360 201 1394
rect 255 1382 288 1399
rect 288 1382 289 1399
rect 255 1365 289 1382
rect 167 1286 201 1320
rect 255 1313 288 1326
rect 288 1313 289 1326
rect 255 1292 289 1313
rect 167 1212 201 1246
rect 255 1244 288 1253
rect 288 1244 289 1253
rect 255 1219 289 1244
rect 255 1175 288 1180
rect 288 1175 289 1180
rect 167 1138 201 1172
rect 255 1146 289 1175
rect 255 1106 288 1107
rect 288 1106 289 1107
rect 167 1064 201 1098
rect 255 1073 289 1106
rect 167 991 201 1025
rect 255 1002 289 1034
rect 255 1000 288 1002
rect 288 1000 289 1002
rect 167 918 201 952
rect 255 933 289 961
rect 255 927 288 933
rect 288 927 289 933
rect 167 845 201 879
rect 255 864 289 888
rect 255 854 288 864
rect 288 854 289 864
rect 167 772 201 806
rect 255 795 289 815
rect 255 781 288 795
rect 288 781 289 795
rect 167 699 201 733
rect 255 726 289 742
rect 255 708 288 726
rect 288 708 289 726
rect 167 626 201 660
rect 255 657 289 670
rect 255 636 288 657
rect 288 636 289 657
rect 255 588 289 598
rect 167 553 201 587
rect 255 564 288 588
rect 288 564 289 588
rect 255 519 289 526
rect 167 480 201 514
rect 255 492 288 519
rect 288 492 289 519
rect 255 450 289 454
rect 167 407 201 441
rect 255 420 288 450
rect 288 420 289 450
rect 255 381 289 382
rect 167 334 201 368
rect 255 348 288 381
rect 288 348 289 381
rect 668 4714 696 4729
rect 696 4714 702 4729
rect 756 4728 790 4762
rect 668 4660 702 4676
rect 539 4634 573 4658
rect 668 4642 696 4660
rect 696 4642 702 4660
rect 756 4655 790 4689
rect 539 4624 546 4634
rect 546 4624 573 4634
rect 668 4591 702 4604
rect 539 4566 573 4583
rect 668 4570 696 4591
rect 696 4570 702 4591
rect 756 4582 790 4616
rect 539 4549 546 4566
rect 546 4549 573 4566
rect 668 4522 702 4532
rect 539 4498 573 4508
rect 668 4498 696 4522
rect 696 4498 702 4522
rect 756 4509 790 4543
rect 539 4474 546 4498
rect 546 4474 573 4498
rect 668 4453 702 4459
rect 539 4430 573 4433
rect 539 4399 546 4430
rect 546 4399 573 4430
rect 668 4425 696 4453
rect 696 4425 702 4453
rect 756 4436 790 4470
rect 668 4384 702 4386
rect 539 4328 546 4357
rect 546 4328 573 4357
rect 668 4352 696 4384
rect 696 4352 702 4384
rect 756 4363 790 4397
rect 539 4323 573 4328
rect 668 4281 696 4313
rect 696 4281 702 4313
rect 756 4290 790 4324
rect 539 4260 546 4281
rect 546 4260 573 4281
rect 668 4279 702 4281
rect 539 4247 573 4260
rect 668 4212 696 4240
rect 696 4212 702 4240
rect 756 4217 790 4251
rect 668 4206 702 4212
rect 539 4192 546 4205
rect 546 4192 573 4205
rect 539 4171 573 4192
rect 668 4143 696 4167
rect 696 4143 702 4167
rect 756 4144 790 4178
rect 668 4133 702 4143
rect 539 4124 546 4129
rect 546 4124 573 4129
rect 539 4095 573 4124
rect 668 4074 696 4094
rect 696 4074 702 4094
rect 668 4060 702 4074
rect 756 4071 790 4105
rect 539 4022 573 4053
rect 539 4019 546 4022
rect 546 4019 573 4022
rect 668 4005 696 4021
rect 696 4005 702 4021
rect 668 3987 702 4005
rect 756 3998 790 4032
rect 539 3954 573 3977
rect 539 3943 546 3954
rect 546 3943 573 3954
rect 668 3936 696 3948
rect 696 3936 702 3948
rect 668 3914 702 3936
rect 756 3925 790 3959
rect 539 3886 573 3901
rect 539 3867 546 3886
rect 546 3867 573 3886
rect 668 3867 696 3875
rect 696 3867 702 3875
rect 668 3841 702 3867
rect 756 3852 790 3886
rect 539 3818 573 3825
rect 539 3791 546 3818
rect 546 3791 573 3818
rect 668 3798 696 3802
rect 696 3798 702 3802
rect 668 3768 702 3798
rect 756 3779 790 3813
rect 668 3695 702 3729
rect 756 3706 790 3740
rect 370 3445 404 3467
rect 370 3433 404 3445
rect 370 3377 404 3393
rect 370 3359 404 3377
rect 370 3309 404 3319
rect 370 3285 404 3309
rect 370 3241 404 3245
rect 370 3211 404 3241
rect 370 3139 404 3171
rect 370 3137 404 3139
rect 370 3071 404 3097
rect 370 3063 404 3071
rect 370 3003 404 3023
rect 370 2989 404 3003
rect 370 2935 404 2950
rect 370 2916 404 2935
rect 370 2867 404 2877
rect 370 2843 404 2867
rect 370 2799 404 2804
rect 370 2770 404 2799
rect 370 1984 404 2016
rect 370 1982 404 1984
rect 370 1916 404 1942
rect 370 1908 404 1916
rect 370 1848 404 1868
rect 370 1834 404 1848
rect 370 1780 404 1794
rect 370 1760 404 1780
rect 370 1712 404 1720
rect 370 1686 404 1712
rect 370 1644 404 1646
rect 370 1612 404 1644
rect 370 1542 404 1572
rect 370 1538 404 1542
rect 370 1464 404 1498
rect 370 1390 404 1424
rect 472 2412 506 2446
rect 472 2340 506 2374
rect 668 3625 702 3656
rect 756 3633 790 3667
rect 668 3622 696 3625
rect 696 3622 702 3625
rect 668 3556 702 3583
rect 756 3559 790 3593
rect 668 3549 696 3556
rect 696 3549 702 3556
rect 668 3487 702 3510
rect 668 3476 696 3487
rect 696 3476 702 3487
rect 756 3485 790 3519
rect 668 3418 702 3437
rect 668 3403 696 3418
rect 696 3403 702 3418
rect 756 3411 790 3445
rect 668 3349 702 3364
rect 668 3330 696 3349
rect 696 3330 702 3349
rect 756 3337 790 3371
rect 668 3280 702 3291
rect 668 3257 696 3280
rect 696 3257 702 3280
rect 756 3263 790 3297
rect 668 3211 702 3218
rect 668 3184 696 3211
rect 696 3184 702 3211
rect 756 3189 790 3223
rect 668 3142 702 3145
rect 668 3111 696 3142
rect 696 3111 702 3142
rect 756 3115 790 3149
rect 668 3039 696 3072
rect 696 3039 702 3072
rect 756 3041 790 3075
rect 668 3038 702 3039
rect 668 2970 696 2999
rect 696 2970 702 2999
rect 668 2965 702 2970
rect 756 2967 790 3001
rect 668 2901 696 2926
rect 696 2901 702 2926
rect 668 2892 702 2901
rect 756 2893 790 2927
rect 668 2832 696 2853
rect 696 2832 702 2853
rect 668 2819 702 2832
rect 756 2819 790 2853
rect 756 2741 790 2775
rect 756 2664 790 2698
rect 756 2587 790 2621
rect 756 2510 790 2544
rect 756 2433 790 2467
rect 756 2356 790 2390
rect 756 2279 790 2313
rect 756 2202 790 2236
rect 756 2124 790 2158
rect 756 2046 790 2080
rect 756 1968 790 2002
rect 668 1900 702 1924
rect 668 1890 696 1900
rect 696 1890 702 1900
rect 756 1890 790 1924
rect 668 1831 702 1851
rect 668 1817 696 1831
rect 696 1817 702 1831
rect 756 1816 790 1850
rect 668 1762 702 1778
rect 668 1744 696 1762
rect 696 1744 702 1762
rect 756 1742 790 1776
rect 668 1693 702 1705
rect 668 1671 696 1693
rect 696 1671 702 1693
rect 756 1668 790 1702
rect 668 1624 702 1632
rect 668 1598 696 1624
rect 696 1598 702 1624
rect 756 1594 790 1628
rect 668 1555 702 1559
rect 668 1525 696 1555
rect 696 1525 702 1555
rect 756 1520 790 1554
rect 668 1452 696 1486
rect 696 1452 702 1486
rect 756 1446 790 1480
rect 370 1316 404 1350
rect 668 1383 696 1413
rect 696 1383 702 1413
rect 668 1379 702 1383
rect 756 1372 790 1406
rect 370 1258 404 1276
rect 370 1242 404 1258
rect 370 1190 404 1202
rect 370 1168 404 1190
rect 370 1122 404 1129
rect 370 1095 404 1122
rect 370 1054 404 1056
rect 370 1022 404 1054
rect 370 952 404 983
rect 370 949 404 952
rect 370 884 404 910
rect 370 876 404 884
rect 370 816 404 837
rect 370 803 404 816
rect 370 748 404 764
rect 370 730 404 748
rect 668 1314 696 1340
rect 696 1314 702 1340
rect 668 1306 702 1314
rect 756 1298 790 1332
rect 668 1245 696 1267
rect 696 1245 702 1267
rect 668 1233 702 1245
rect 756 1224 790 1258
rect 668 1176 696 1194
rect 696 1176 702 1194
rect 668 1160 702 1176
rect 756 1150 790 1184
rect 668 1107 696 1121
rect 696 1107 702 1121
rect 668 1087 702 1107
rect 756 1076 790 1110
rect 668 1038 696 1048
rect 696 1038 702 1048
rect 668 1014 702 1038
rect 756 1002 790 1036
rect 668 969 696 975
rect 696 969 702 975
rect 668 941 702 969
rect 756 928 790 962
rect 668 900 696 902
rect 696 900 702 902
rect 668 868 702 900
rect 756 854 790 888
rect 668 796 702 828
rect 668 794 696 796
rect 696 794 702 796
rect 756 780 790 814
rect 668 727 702 754
rect 668 720 696 727
rect 696 720 702 727
rect 756 706 790 740
rect 668 658 702 680
rect 668 646 696 658
rect 696 646 702 658
rect 756 632 790 666
rect 668 589 702 606
rect 668 572 696 589
rect 696 572 702 589
rect 756 558 790 592
rect 668 520 702 532
rect 668 498 696 520
rect 696 498 702 520
rect 756 484 790 518
rect 668 451 702 458
rect 668 424 696 451
rect 696 424 702 451
rect 756 410 790 444
rect 668 382 702 384
rect 668 350 696 382
rect 696 350 702 382
rect 756 335 790 369
rect 167 261 201 295
rect 255 278 288 310
rect 288 278 289 310
rect 255 276 289 278
rect 338 288 372 310
rect 421 288 455 310
rect 504 288 538 310
rect 586 288 620 310
rect 668 288 702 310
rect 338 276 352 288
rect 352 276 372 288
rect 421 276 423 288
rect 423 276 455 288
rect 504 276 528 288
rect 528 276 538 288
rect 586 276 600 288
rect 600 276 620 288
rect 668 276 672 288
rect 672 276 702 288
rect 756 260 790 294
rect 239 188 273 222
rect 313 188 347 222
rect 387 188 421 222
rect 461 188 495 222
rect 535 188 569 222
rect 609 188 643 222
rect 683 188 717 222
rect -44 81 -10 115
rect 59 68 92 101
rect 92 68 93 101
rect 134 68 161 101
rect 161 68 168 101
rect 209 68 230 101
rect 230 68 243 101
rect 284 68 300 101
rect 300 68 318 101
rect 359 68 370 101
rect 370 68 393 101
rect 434 68 440 101
rect 440 68 468 101
rect 509 68 510 101
rect 510 68 543 101
rect 584 68 614 101
rect 614 68 618 101
rect 659 68 684 101
rect 684 68 693 101
rect 734 68 754 101
rect 754 68 768 101
rect 808 68 824 101
rect 824 68 842 101
rect 59 67 93 68
rect 134 67 168 68
rect 209 67 243 68
rect 284 67 318 68
rect 359 67 393 68
rect 434 67 468 68
rect 509 67 543 68
rect 584 67 618 68
rect 659 67 693 68
rect 734 67 768 68
rect 808 67 842 68
rect -44 7 -10 41
<< metal1 >>
rect -26 12129 92 12141
rect -26 12095 -20 12129
rect 14 12095 52 12129
rect 86 12095 92 12129
rect -26 12055 92 12095
rect -26 12021 -20 12055
rect 14 12021 52 12055
rect 86 12021 92 12055
rect -26 11981 92 12021
rect 151 12044 776 12050
rect 151 12010 163 12044
rect 197 12010 246 12044
rect 280 12010 329 12044
rect 363 12010 412 12044
rect 446 12010 496 12044
rect 530 12010 580 12044
rect 614 12010 664 12044
rect 698 12010 776 12044
rect 151 12004 776 12010
rect -26 11947 -20 11981
rect 14 11947 52 11981
rect 86 11947 92 11981
rect -26 11907 92 11947
rect -26 11873 -20 11907
rect 14 11873 52 11907
rect 86 11873 92 11907
rect -26 11833 92 11873
rect -26 11799 -20 11833
rect 14 11799 52 11833
rect 86 11799 92 11833
rect -26 11759 92 11799
rect -26 11725 -20 11759
rect 14 11725 52 11759
rect 86 11725 92 11759
rect -26 11685 92 11725
rect -26 11651 -20 11685
rect 14 11651 52 11685
rect 86 11651 92 11685
rect -26 11611 92 11651
rect -26 11577 -20 11611
rect 14 11577 52 11611
rect 86 11577 92 11611
rect -26 11537 92 11577
rect -26 11503 -20 11537
rect 14 11503 52 11537
rect 86 11503 92 11537
rect -26 11463 92 11503
rect -26 11429 -20 11463
rect 14 11429 52 11463
rect 86 11429 92 11463
rect -26 11389 92 11429
rect -26 11355 -20 11389
rect 14 11355 52 11389
rect 86 11355 92 11389
rect -26 11315 92 11355
rect -26 11281 -20 11315
rect 14 11281 52 11315
rect 86 11281 92 11315
rect -26 11241 92 11281
rect -26 11207 -20 11241
rect 14 11207 52 11241
rect 86 11207 92 11241
rect -26 11167 92 11207
rect -26 11133 -20 11167
rect 14 11133 52 11167
rect 86 11133 92 11167
rect -26 11093 92 11133
rect -26 11059 -20 11093
rect 14 11059 52 11093
rect 86 11059 92 11093
rect -26 11019 92 11059
rect -26 10985 -20 11019
rect 14 10985 52 11019
rect 86 10985 92 11019
rect -26 10945 92 10985
rect -26 10911 -20 10945
rect 14 10911 52 10945
rect 86 10911 92 10945
rect -26 10871 92 10911
rect -26 10837 -20 10871
rect 14 10837 52 10871
rect 86 10837 92 10871
rect -26 10797 92 10837
rect -26 10763 -20 10797
rect 14 10763 52 10797
rect 86 10763 92 10797
rect -26 10723 92 10763
rect -26 10689 -20 10723
rect 14 10689 52 10723
rect 86 10689 92 10723
rect -26 10649 92 10689
rect -26 10615 -20 10649
rect 14 10615 52 10649
rect 86 10615 92 10649
rect -26 10575 92 10615
rect -26 10541 -20 10575
rect 14 10541 52 10575
rect 86 10541 92 10575
rect -26 10502 92 10541
rect -26 10468 -20 10502
rect 14 10468 52 10502
rect 86 10468 92 10502
rect -26 10429 92 10468
rect -26 10395 -20 10429
rect 14 10395 52 10429
rect 86 10395 92 10429
rect -26 10356 92 10395
rect -26 10322 -20 10356
rect 14 10322 52 10356
rect 86 10322 92 10356
rect -26 10283 92 10322
rect -26 10249 -20 10283
rect 14 10249 52 10283
rect 86 10249 92 10283
rect -26 10210 92 10249
rect -26 10176 -20 10210
rect 14 10176 52 10210
rect 86 10176 92 10210
rect -26 10137 92 10176
rect -26 10103 -20 10137
rect 14 10103 52 10137
rect 86 10103 92 10137
rect -26 10064 92 10103
rect -26 10030 -20 10064
rect 14 10030 52 10064
rect 86 10030 92 10064
rect -26 9991 92 10030
rect -26 9957 -20 9991
rect 14 9957 52 9991
rect 86 9957 92 9991
rect -26 9918 92 9957
rect -26 9884 -20 9918
rect 14 9884 52 9918
rect 86 9884 92 9918
rect -26 9845 92 9884
rect -26 9811 -20 9845
rect 14 9811 52 9845
rect 86 9811 92 9845
rect 152 11972 776 12004
rect 152 11959 736 11972
rect 152 11925 230 11959
rect 264 11925 302 11959
rect 336 11925 374 11959
rect 408 11925 446 11959
rect 480 11925 518 11959
rect 552 11925 590 11959
rect 624 11938 736 11959
rect 770 11938 776 11972
rect 624 11925 776 11938
rect 152 11900 776 11925
rect 152 11887 736 11900
rect 152 11853 158 11887
rect 192 11853 662 11887
rect 696 11866 736 11887
rect 770 11866 776 11900
rect 696 11853 776 11866
rect 152 11828 776 11853
rect 152 11815 736 11828
rect 152 11811 662 11815
rect 152 11777 158 11811
rect 192 11781 662 11811
rect 696 11794 736 11815
rect 770 11794 776 11828
rect 696 11781 776 11794
rect 192 11777 776 11781
rect 152 11756 776 11777
rect 152 11743 736 11756
rect 152 11735 662 11743
rect 152 11701 158 11735
rect 192 11709 662 11735
rect 696 11722 736 11743
rect 770 11722 776 11756
rect 696 11709 776 11722
rect 192 11701 776 11709
rect 152 11684 776 11701
rect 152 11671 736 11684
rect 152 11659 662 11671
rect 152 11625 158 11659
rect 192 11637 662 11659
rect 696 11650 736 11671
rect 770 11650 776 11684
rect 696 11637 776 11650
rect 192 11625 776 11637
rect 152 11612 776 11625
rect 152 11599 736 11612
rect 152 11583 662 11599
rect 152 11549 158 11583
rect 192 11565 662 11583
rect 696 11578 736 11599
rect 770 11578 776 11612
rect 696 11565 776 11578
rect 192 11549 776 11565
rect 152 11540 776 11549
rect 152 11527 736 11540
rect 152 11507 662 11527
rect 152 11473 158 11507
rect 192 11493 662 11507
rect 696 11506 736 11527
rect 770 11506 776 11540
rect 696 11493 776 11506
rect 192 11473 776 11493
rect 152 11468 776 11473
rect 152 11455 736 11468
rect 152 11431 662 11455
rect 152 11397 158 11431
rect 192 11421 662 11431
rect 696 11434 736 11455
rect 770 11434 776 11468
rect 696 11421 776 11434
rect 192 11397 776 11421
rect 152 11396 776 11397
rect 152 11383 736 11396
rect 152 11355 662 11383
rect 152 11321 158 11355
rect 192 11349 662 11355
rect 696 11362 736 11383
rect 770 11362 776 11396
rect 696 11349 776 11362
rect 192 11324 776 11349
rect 192 11321 736 11324
rect 152 11311 736 11321
rect 152 11279 662 11311
rect 152 11245 158 11279
rect 192 11277 662 11279
rect 696 11290 736 11311
rect 770 11290 776 11324
rect 696 11277 776 11290
rect 192 11252 776 11277
rect 192 11245 736 11252
rect 152 11239 736 11245
rect 152 11205 662 11239
rect 696 11218 736 11239
rect 770 11218 776 11252
rect 696 11205 776 11218
rect 152 11203 776 11205
rect 152 11169 158 11203
rect 192 11180 776 11203
rect 192 11169 736 11180
rect 152 11167 736 11169
rect 152 11133 662 11167
rect 696 11146 736 11167
rect 770 11146 776 11180
rect 696 11133 776 11146
rect 152 11127 776 11133
rect 152 11093 158 11127
rect 192 11108 776 11127
rect 192 11095 736 11108
rect 192 11093 662 11095
rect 152 11061 662 11093
rect 696 11074 736 11095
rect 770 11074 776 11108
rect 696 11061 776 11074
rect 152 11051 776 11061
rect 152 11017 158 11051
rect 192 11036 776 11051
rect 192 11023 736 11036
rect 192 11017 662 11023
rect 152 10989 662 11017
rect 696 11002 736 11023
rect 770 11002 776 11036
rect 696 10989 776 11002
rect 152 10975 776 10989
rect 152 10941 158 10975
rect 192 10964 776 10975
rect 192 10951 736 10964
rect 192 10941 662 10951
rect 152 10917 662 10941
rect 696 10930 736 10951
rect 770 10930 776 10964
rect 696 10917 776 10930
rect 152 10899 776 10917
rect 152 10865 158 10899
rect 192 10892 776 10899
rect 192 10879 736 10892
rect 192 10865 662 10879
rect 152 10845 662 10865
rect 696 10858 736 10879
rect 770 10858 776 10892
rect 696 10845 776 10858
rect 152 10823 776 10845
rect 152 10789 158 10823
rect 192 10820 776 10823
rect 192 10807 736 10820
rect 192 10789 662 10807
rect 152 10773 662 10789
rect 696 10786 736 10807
rect 770 10786 776 10820
rect 696 10773 776 10786
rect 152 10748 776 10773
rect 152 10747 736 10748
rect 152 10713 158 10747
rect 192 10735 736 10747
rect 192 10713 662 10735
rect 152 10701 662 10713
rect 696 10714 736 10735
rect 770 10714 776 10748
rect 696 10701 776 10714
rect 152 10676 776 10701
rect 152 10672 736 10676
rect 152 10638 158 10672
rect 192 10663 736 10672
rect 192 10645 662 10663
rect 192 10638 318 10645
rect 152 10597 318 10638
rect 152 10563 158 10597
rect 192 10563 318 10597
rect 152 10522 318 10563
rect 152 10488 158 10522
rect 192 10488 318 10522
rect 152 10439 318 10488
rect 152 10405 158 10439
rect 192 10405 278 10439
rect 312 10405 318 10439
rect 152 10360 318 10405
rect 152 10326 158 10360
rect 192 10326 278 10360
rect 312 10326 318 10360
rect 152 10292 318 10326
rect 152 10240 154 10292
rect 206 10240 258 10292
rect 310 10281 318 10292
rect 312 10247 318 10281
rect 310 10240 318 10247
rect 152 10202 318 10240
rect 152 10188 158 10202
rect 192 10188 278 10202
rect 152 10136 154 10188
rect 206 10136 258 10188
rect 312 10168 318 10202
rect 310 10136 318 10168
rect 152 10123 318 10136
rect 152 10089 158 10123
rect 192 10089 278 10123
rect 312 10089 318 10123
rect 152 10083 318 10089
rect 152 10031 154 10083
rect 206 10031 258 10083
rect 310 10043 318 10083
rect 152 10009 158 10031
rect 192 10009 278 10031
rect 312 10009 318 10043
rect 152 9978 318 10009
rect 152 9926 154 9978
rect 206 9926 258 9978
rect 310 9963 318 9978
rect 312 9929 318 9963
rect 310 9926 318 9929
rect 152 9883 318 9926
rect 152 9873 158 9883
rect 192 9873 278 9883
rect 152 9837 154 9873
rect -26 9772 92 9811
rect -26 9738 -20 9772
rect 14 9738 52 9772
rect 86 9738 92 9772
rect -26 9699 92 9738
rect 206 9821 258 9873
rect 312 9849 318 9883
rect 310 9837 318 9849
rect 656 10629 662 10645
rect 696 10642 736 10663
rect 770 10642 776 10676
rect 696 10629 776 10642
rect 656 10604 776 10629
rect 656 10591 736 10604
rect 656 10557 662 10591
rect 696 10570 736 10591
rect 770 10570 776 10604
rect 696 10557 776 10570
rect 656 10532 776 10557
rect 656 10519 736 10532
rect 656 10485 662 10519
rect 696 10498 736 10519
rect 770 10498 776 10532
rect 696 10485 776 10498
rect 656 10460 776 10485
rect 656 10447 736 10460
rect 656 10413 662 10447
rect 696 10426 736 10447
rect 770 10426 776 10460
rect 696 10413 776 10426
rect 656 10388 776 10413
rect 656 10375 736 10388
rect 656 10341 662 10375
rect 696 10354 736 10375
rect 770 10354 776 10388
rect 696 10341 776 10354
rect 656 10316 776 10341
rect 656 10303 736 10316
rect 656 10269 662 10303
rect 696 10282 736 10303
rect 770 10282 776 10316
rect 696 10269 776 10282
rect 656 10244 776 10269
rect 656 10231 736 10244
rect 656 10197 662 10231
rect 696 10210 736 10231
rect 770 10210 776 10244
rect 696 10197 776 10210
rect 656 10172 776 10197
rect 656 10159 736 10172
rect 656 10125 662 10159
rect 696 10138 736 10159
rect 770 10138 776 10172
rect 696 10125 776 10138
rect 656 10100 776 10125
rect 656 10087 736 10100
rect 656 10053 662 10087
rect 696 10066 736 10087
rect 770 10066 776 10100
rect 696 10053 776 10066
rect 656 10028 776 10053
rect 656 10015 736 10028
rect 656 9981 662 10015
rect 696 9994 736 10015
rect 770 9994 776 10028
rect 696 9981 776 9994
rect 656 9956 776 9981
rect 656 9943 736 9956
rect 656 9909 662 9943
rect 696 9922 736 9943
rect 770 9922 776 9956
rect 696 9909 776 9922
rect 656 9884 776 9909
rect 656 9871 736 9884
rect 656 9837 662 9871
rect 696 9850 736 9871
rect 770 9850 776 9884
rect 696 9837 776 9850
rect 154 9768 310 9821
rect 206 9716 258 9768
rect 154 9710 310 9716
rect 656 9812 776 9837
rect 656 9799 736 9812
rect 656 9765 662 9799
rect 696 9778 736 9799
rect 770 9778 776 9812
rect 696 9765 776 9778
rect 656 9740 776 9765
rect 656 9727 736 9740
rect -26 9665 -20 9699
rect 14 9665 52 9699
rect 86 9665 92 9699
rect -26 9626 92 9665
rect -26 9592 -20 9626
rect 14 9592 52 9626
rect 86 9592 92 9626
rect -26 9553 92 9592
rect -26 9519 -20 9553
rect 14 9519 52 9553
rect 86 9519 92 9553
rect -26 9480 92 9519
rect -26 9446 -20 9480
rect 14 9446 52 9480
rect 86 9446 92 9480
rect -26 9434 92 9446
rect 656 9693 662 9727
rect 696 9706 736 9727
rect 770 9706 776 9740
rect 696 9693 776 9706
rect 656 9668 776 9693
rect 656 9655 736 9668
rect 656 9621 662 9655
rect 696 9634 736 9655
rect 770 9634 776 9668
rect 696 9621 776 9634
rect 656 9596 776 9621
rect 656 9583 736 9596
rect 656 9549 662 9583
rect 696 9562 736 9583
rect 770 9562 776 9596
rect 696 9549 776 9562
rect 656 9524 776 9549
rect 656 9511 736 9524
rect 656 9477 662 9511
rect 696 9490 736 9511
rect 770 9490 776 9524
rect 696 9477 776 9490
rect 656 9452 776 9477
rect 656 9439 736 9452
rect 656 9405 662 9439
rect 696 9418 736 9439
rect 770 9418 776 9452
rect 696 9405 776 9418
rect 656 9380 776 9405
rect 656 9367 736 9380
rect 656 9333 662 9367
rect 696 9346 736 9367
rect 770 9346 776 9380
rect 696 9333 776 9346
rect 656 9308 776 9333
rect 656 9294 736 9308
rect 656 9260 662 9294
rect 696 9274 736 9294
rect 770 9274 776 9308
rect 696 9260 776 9274
rect 656 9236 776 9260
rect 656 9221 736 9236
rect 656 9187 662 9221
rect 696 9202 736 9221
rect 770 9202 776 9236
rect 696 9187 776 9202
rect -26 9163 92 9175
rect -26 9129 -20 9163
rect 14 9129 52 9163
rect 86 9129 92 9163
rect -26 9088 92 9129
rect -26 9054 -20 9088
rect 14 9054 52 9088
rect 86 9054 92 9088
rect -26 9013 92 9054
rect -26 8979 -20 9013
rect 14 8979 52 9013
rect 86 8979 92 9013
rect -26 8938 92 8979
rect -26 8904 -20 8938
rect 14 8904 52 8938
rect 86 8904 92 8938
rect -26 8863 92 8904
rect -26 8829 -20 8863
rect 14 8829 52 8863
rect 86 8829 92 8863
rect -26 8788 92 8829
rect -26 8754 -20 8788
rect 14 8754 52 8788
rect 86 8754 92 8788
rect -26 8713 92 8754
rect -26 8679 -20 8713
rect 14 8679 52 8713
rect 86 8679 92 8713
rect -26 8638 92 8679
rect -26 8604 -20 8638
rect 14 8604 52 8638
rect 86 8604 92 8638
rect 656 9164 776 9187
rect 656 9148 736 9164
rect 656 9114 662 9148
rect 696 9130 736 9148
rect 770 9130 776 9164
rect 696 9114 776 9130
rect 656 9092 776 9114
rect 656 9075 736 9092
rect 656 9041 662 9075
rect 696 9058 736 9075
rect 770 9058 776 9092
rect 696 9041 776 9058
rect 656 9020 776 9041
rect 656 9002 736 9020
rect 656 8968 662 9002
rect 696 8986 736 9002
rect 770 8986 776 9020
rect 696 8968 776 8986
rect 656 8948 776 8968
rect 656 8929 736 8948
rect 656 8895 662 8929
rect 696 8914 736 8929
rect 770 8914 776 8948
rect 696 8895 776 8914
rect 656 8876 776 8895
rect 656 8856 736 8876
rect 656 8822 662 8856
rect 696 8842 736 8856
rect 770 8842 776 8876
rect 696 8822 776 8842
rect 656 8804 776 8822
rect 656 8783 736 8804
rect 656 8749 662 8783
rect 696 8770 736 8783
rect 770 8770 776 8804
rect 696 8749 776 8770
rect 656 8732 776 8749
rect 656 8710 736 8732
rect 656 8676 662 8710
rect 696 8698 736 8710
rect 770 8698 776 8732
rect 696 8676 776 8698
rect 656 8660 776 8676
rect 656 8637 736 8660
rect -26 8563 92 8604
rect -26 8529 -20 8563
rect 14 8529 52 8563
rect 86 8529 92 8563
rect -26 8488 92 8529
rect -26 8454 -20 8488
rect 14 8454 52 8488
rect 86 8454 92 8488
rect -26 8413 92 8454
rect -26 8379 -20 8413
rect 14 8379 52 8413
rect 86 8379 92 8413
rect -26 8338 92 8379
rect -26 8304 -20 8338
rect 14 8304 52 8338
rect 86 8304 92 8338
rect -26 8263 92 8304
rect -26 8229 -20 8263
rect 14 8229 52 8263
rect 86 8229 92 8263
rect -26 8188 92 8229
rect -26 8154 -20 8188
rect 14 8154 52 8188
rect 86 8154 92 8188
rect -26 8113 92 8154
rect -26 8079 -20 8113
rect 14 8079 52 8113
rect 86 8079 92 8113
rect -26 8038 92 8079
rect -26 8004 -20 8038
rect 14 8004 52 8038
rect 86 8004 92 8038
rect 152 8621 318 8633
rect 152 8587 158 8621
rect 192 8587 278 8621
rect 312 8587 318 8621
rect 152 8542 318 8587
rect 152 8508 158 8542
rect 192 8508 278 8542
rect 312 8508 318 8542
rect 152 8477 318 8508
rect 152 8425 154 8477
rect 206 8425 258 8477
rect 310 8463 318 8477
rect 312 8429 318 8463
rect 310 8425 318 8429
rect 152 8412 318 8425
rect 152 8360 154 8412
rect 206 8360 258 8412
rect 310 8384 318 8412
rect 152 8350 158 8360
rect 192 8350 278 8360
rect 312 8350 318 8384
rect 152 8347 318 8350
rect 152 8295 154 8347
rect 206 8295 258 8347
rect 310 8305 318 8347
rect 152 8282 158 8295
rect 192 8282 278 8295
rect 152 8230 154 8282
rect 206 8230 258 8282
rect 312 8271 318 8305
rect 310 8230 318 8271
rect 152 8225 318 8230
rect 152 8217 158 8225
rect 192 8217 278 8225
rect 152 8165 154 8217
rect 206 8165 258 8217
rect 312 8191 318 8225
rect 310 8165 318 8191
rect 152 8151 318 8165
rect 152 8099 154 8151
rect 206 8099 258 8151
rect 310 8145 318 8151
rect 312 8111 318 8145
rect 310 8099 318 8111
rect 152 8085 318 8099
rect 152 8033 154 8085
rect 206 8033 258 8085
rect 310 8065 318 8085
rect 152 8031 158 8033
rect 192 8031 278 8033
rect 312 8031 318 8065
rect 152 8019 318 8031
rect 656 8603 662 8637
rect 696 8626 736 8637
rect 770 8626 776 8660
rect 696 8603 776 8626
rect 656 8588 776 8603
rect 656 8564 736 8588
rect 656 8530 662 8564
rect 696 8554 736 8564
rect 770 8554 776 8588
rect 696 8530 776 8554
rect 656 8516 776 8530
rect 656 8491 736 8516
rect 656 8457 662 8491
rect 696 8482 736 8491
rect 770 8482 776 8516
rect 696 8457 776 8482
rect 656 8444 776 8457
rect 656 8418 736 8444
rect 656 8384 662 8418
rect 696 8410 736 8418
rect 770 8410 776 8444
rect 696 8384 776 8410
rect 656 8372 776 8384
rect 656 8345 736 8372
rect 656 8311 662 8345
rect 696 8338 736 8345
rect 770 8338 776 8372
rect 696 8311 776 8338
rect 656 8300 776 8311
rect 656 8272 736 8300
rect 656 8238 662 8272
rect 696 8266 736 8272
rect 770 8266 776 8300
rect 696 8238 776 8266
rect 656 8228 776 8238
rect 656 8199 736 8228
rect 656 8165 662 8199
rect 696 8194 736 8199
rect 770 8194 776 8228
rect 696 8165 776 8194
rect 656 8156 776 8165
rect 656 8126 736 8156
rect 656 8092 662 8126
rect 696 8122 736 8126
rect 770 8122 776 8156
rect 696 8092 776 8122
rect 656 8084 776 8092
rect 656 8053 736 8084
rect 656 8019 662 8053
rect 696 8050 736 8053
rect 770 8050 776 8084
rect 696 8019 776 8050
rect -26 7963 92 8004
rect -26 7929 -20 7963
rect 14 7929 52 7963
rect 86 7929 92 7963
rect -26 7889 92 7929
rect 206 7967 258 8019
rect 154 7953 310 7967
rect 206 7901 258 7953
rect 154 7895 310 7901
rect 656 8012 776 8019
rect 656 7980 736 8012
rect 656 7946 662 7980
rect 696 7978 736 7980
rect 770 7978 776 8012
rect 696 7946 776 7978
rect 656 7940 776 7946
rect 656 7907 736 7940
rect -26 7855 -20 7889
rect 14 7855 52 7889
rect 86 7855 92 7889
rect -26 7815 92 7855
rect -26 7781 -20 7815
rect 14 7781 52 7815
rect 86 7781 92 7815
rect -26 7741 92 7781
rect -26 7707 -20 7741
rect 14 7707 52 7741
rect 86 7707 92 7741
rect -26 7667 92 7707
rect -26 7640 -20 7667
rect -191 7633 -20 7640
rect 14 7633 52 7667
rect 86 7633 92 7667
rect -191 7593 92 7633
rect -191 7559 -20 7593
rect 14 7559 52 7593
rect 86 7559 92 7593
rect -191 7547 92 7559
rect 656 7873 662 7907
rect 696 7906 736 7907
rect 770 7906 776 7940
rect 696 7873 776 7906
rect 656 7868 776 7873
rect 656 7834 736 7868
rect 770 7834 776 7868
rect 656 7800 662 7834
rect 696 7800 776 7834
rect 656 7796 776 7800
rect 656 7762 736 7796
rect 770 7762 776 7796
rect 656 7761 776 7762
rect 656 7727 662 7761
rect 696 7727 776 7761
rect 656 7724 776 7727
rect 656 7690 736 7724
rect 770 7690 776 7724
rect 656 7688 776 7690
rect 656 7654 662 7688
rect 696 7654 776 7688
rect 656 7652 776 7654
rect 656 7618 736 7652
rect 770 7618 776 7652
rect 656 7615 776 7618
rect 656 7581 662 7615
rect 696 7581 776 7615
rect 656 7580 776 7581
rect -191 7280 -142 7547
rect 656 7546 736 7580
rect 770 7546 776 7580
rect 656 7542 776 7546
rect 656 7508 662 7542
rect 696 7508 776 7542
rect 656 7474 736 7508
rect 770 7474 776 7508
rect 656 7469 776 7474
rect 656 7435 662 7469
rect 696 7436 776 7469
rect 696 7435 736 7436
rect 656 7402 736 7435
rect 770 7402 776 7436
rect 656 7396 776 7402
rect 656 7362 662 7396
rect 696 7364 776 7396
rect 696 7362 736 7364
rect 656 7330 736 7362
rect 770 7330 776 7364
rect 656 7323 776 7330
rect 656 7289 662 7323
rect 696 7292 776 7323
rect 696 7289 736 7292
rect -191 7268 92 7280
rect -191 7234 -20 7268
rect 14 7234 52 7268
rect 86 7234 92 7268
rect -191 7194 92 7234
rect -191 7190 -20 7194
rect -26 7160 -20 7190
rect 14 7160 52 7194
rect 86 7160 92 7194
rect -26 7120 92 7160
rect -26 7086 -20 7120
rect 14 7086 52 7120
rect 86 7086 92 7120
rect -26 7046 92 7086
rect -26 7012 -20 7046
rect 14 7012 52 7046
rect 86 7012 92 7046
rect -26 6972 92 7012
rect -26 6938 -20 6972
rect 14 6938 52 6972
rect 86 6938 92 6972
rect -26 6898 92 6938
rect -26 6864 -20 6898
rect 14 6864 52 6898
rect 86 6864 92 6898
rect -26 6824 92 6864
rect -26 6790 -20 6824
rect 14 6790 52 6824
rect 86 6790 92 6824
rect -26 6750 92 6790
rect -26 6716 -20 6750
rect 14 6716 52 6750
rect 86 6716 92 6750
rect -26 6676 92 6716
rect -26 6642 -20 6676
rect 14 6642 52 6676
rect 86 6642 92 6676
rect -26 6602 92 6642
rect -26 6568 -20 6602
rect 14 6568 52 6602
rect 86 6568 92 6602
rect -26 6528 92 6568
rect -26 6494 -20 6528
rect 14 6494 52 6528
rect 86 6494 92 6528
rect -26 6454 92 6494
rect -26 6420 -20 6454
rect 14 6420 52 6454
rect 86 6420 92 6454
rect -26 6380 92 6420
rect -26 6346 -20 6380
rect 14 6346 52 6380
rect 86 6346 92 6380
rect -26 6306 92 6346
rect -26 6272 -20 6306
rect 14 6272 52 6306
rect 86 6272 92 6306
rect -26 6233 92 6272
rect -26 6199 -20 6233
rect 14 6199 52 6233
rect 86 6199 92 6233
rect -26 6160 92 6199
rect -26 6126 -20 6160
rect 14 6126 52 6160
rect 86 6126 92 6160
rect -26 6087 92 6126
rect -26 6053 -20 6087
rect 14 6053 52 6087
rect 86 6053 92 6087
rect -26 6014 92 6053
rect -26 5980 -20 6014
rect 14 5980 52 6014
rect 86 5980 92 6014
rect -26 5941 92 5980
rect -26 5907 -20 5941
rect 14 5907 52 5941
rect 86 5907 92 5941
rect -26 5868 92 5907
rect -26 5834 -20 5868
rect 14 5834 52 5868
rect 86 5834 92 5868
rect -26 5795 92 5834
rect -26 5761 -20 5795
rect 14 5761 52 5795
rect 86 5761 92 5795
rect -26 5722 92 5761
rect -26 5688 -20 5722
rect 14 5688 52 5722
rect 86 5688 92 5722
rect -26 5649 92 5688
rect -26 5615 -20 5649
rect 14 5615 52 5649
rect 86 5615 92 5649
rect -26 5576 92 5615
rect -26 5542 -20 5576
rect 14 5542 52 5576
rect 86 5542 92 5576
rect -26 5503 92 5542
rect -26 5469 -20 5503
rect 14 5469 52 5503
rect 86 5469 92 5503
rect -26 5430 92 5469
rect -26 5396 -20 5430
rect 14 5396 52 5430
rect 86 5396 92 5430
rect -26 5357 92 5396
rect -26 5323 -20 5357
rect 14 5323 52 5357
rect 86 5323 92 5357
rect -26 5284 92 5323
rect -26 5250 -20 5284
rect 14 5250 52 5284
rect 86 5250 92 5284
rect -26 5211 92 5250
rect -26 5177 -20 5211
rect 14 5177 52 5211
rect 86 5177 92 5211
rect -26 5138 92 5177
rect -26 5104 -20 5138
rect 14 5104 52 5138
rect 86 5104 92 5138
rect -26 5065 92 5104
rect 153 7273 223 7285
rect 153 7239 171 7273
rect 205 7239 223 7273
rect 153 7199 223 7239
rect 153 7165 171 7199
rect 205 7165 223 7199
rect 153 7125 223 7165
rect 153 7091 171 7125
rect 205 7091 223 7125
rect 153 7087 223 7091
rect 153 7035 162 7087
rect 214 7035 223 7087
rect 153 7022 171 7035
rect 205 7022 223 7035
rect 153 6970 162 7022
rect 214 6970 223 7022
rect 153 6957 171 6970
rect 205 6957 223 6970
rect 153 6905 162 6957
rect 214 6905 223 6957
rect 153 6892 171 6905
rect 205 6892 223 6905
rect 153 6840 162 6892
rect 214 6840 223 6892
rect 153 6833 223 6840
rect 153 6826 171 6833
rect 205 6826 223 6833
rect 153 6774 162 6826
rect 214 6774 223 6826
rect 153 6760 223 6774
rect 153 6708 162 6760
rect 214 6708 223 6760
rect 153 6694 223 6708
rect 153 6642 162 6694
rect 214 6642 223 6694
rect 153 6628 223 6642
rect 153 6576 162 6628
rect 214 6576 223 6628
rect 153 6562 223 6576
rect 153 6510 162 6562
rect 214 6510 223 6562
rect 153 6507 171 6510
rect 205 6507 223 6510
rect 153 6496 223 6507
rect 153 6444 162 6496
rect 214 6444 223 6496
rect 153 6434 171 6444
rect 205 6434 223 6444
rect 153 6430 223 6434
rect 153 6378 162 6430
rect 214 6378 223 6430
rect 153 6364 171 6378
rect 205 6364 223 6378
rect 153 6312 162 6364
rect 214 6312 223 6364
rect 153 6298 171 6312
rect 205 6298 223 6312
rect 153 6246 162 6298
rect 214 6246 223 6298
rect 153 6232 171 6246
rect 205 6232 223 6246
rect 153 6180 162 6232
rect 214 6180 223 6232
rect 153 6176 223 6180
rect 153 6166 171 6176
rect 205 6166 223 6176
rect 153 6114 162 6166
rect 214 6121 223 6166
rect 656 7258 736 7289
rect 770 7258 776 7292
rect 656 7250 776 7258
rect 656 7216 662 7250
rect 696 7220 776 7250
rect 696 7216 736 7220
rect 656 7186 736 7216
rect 770 7186 776 7220
rect 656 7177 776 7186
rect 656 7143 662 7177
rect 696 7148 776 7177
rect 696 7143 736 7148
rect 656 7114 736 7143
rect 770 7114 776 7148
rect 656 7104 776 7114
rect 656 7070 662 7104
rect 696 7076 776 7104
rect 696 7070 736 7076
rect 656 7042 736 7070
rect 770 7042 776 7076
rect 656 7031 776 7042
rect 656 6997 662 7031
rect 696 7004 776 7031
rect 696 6997 736 7004
rect 656 6970 736 6997
rect 770 6970 776 7004
rect 656 6958 776 6970
rect 656 6924 662 6958
rect 696 6932 776 6958
rect 696 6924 736 6932
rect 656 6898 736 6924
rect 770 6898 776 6932
rect 656 6885 776 6898
rect 656 6851 662 6885
rect 696 6860 776 6885
rect 696 6851 736 6860
rect 656 6826 736 6851
rect 770 6826 776 6860
rect 656 6812 776 6826
rect 656 6778 662 6812
rect 696 6788 776 6812
rect 696 6778 736 6788
rect 656 6754 736 6778
rect 770 6754 776 6788
rect 656 6739 776 6754
rect 656 6705 662 6739
rect 696 6716 776 6739
rect 696 6705 736 6716
rect 656 6682 736 6705
rect 770 6682 776 6716
rect 656 6666 776 6682
rect 656 6632 662 6666
rect 696 6644 776 6666
rect 696 6632 736 6644
rect 656 6610 736 6632
rect 770 6610 776 6644
rect 656 6593 776 6610
rect 656 6559 662 6593
rect 696 6572 776 6593
rect 696 6559 736 6572
rect 656 6538 736 6559
rect 770 6538 776 6572
rect 656 6520 776 6538
rect 656 6486 662 6520
rect 696 6500 776 6520
rect 696 6486 736 6500
rect 656 6466 736 6486
rect 770 6466 776 6500
rect 656 6447 776 6466
rect 656 6413 662 6447
rect 696 6428 776 6447
rect 696 6413 736 6428
rect 656 6394 736 6413
rect 770 6394 776 6428
rect 656 6374 776 6394
rect 656 6340 662 6374
rect 696 6356 776 6374
rect 696 6340 736 6356
rect 656 6322 736 6340
rect 770 6322 776 6356
rect 656 6301 776 6322
rect 656 6267 662 6301
rect 696 6284 776 6301
rect 696 6267 736 6284
rect 656 6250 736 6267
rect 770 6250 776 6284
rect 656 6228 776 6250
rect 656 6194 662 6228
rect 696 6212 776 6228
rect 696 6194 736 6212
rect 656 6178 736 6194
rect 770 6178 776 6212
rect 656 6155 776 6178
tri 223 6121 234 6132 sw
rect 656 6121 662 6155
rect 696 6140 776 6155
rect 696 6121 736 6140
rect 214 6114 234 6121
rect 153 6106 234 6114
tri 234 6106 249 6121 sw
rect 656 6106 736 6121
rect 770 6106 776 6140
rect 153 6103 249 6106
rect 153 6100 171 6103
rect 205 6100 249 6103
rect 153 6048 162 6100
rect 214 6082 249 6100
tri 249 6082 273 6106 sw
rect 656 6082 776 6106
rect 214 6077 273 6082
tri 273 6077 278 6082 sw
rect 656 6077 662 6082
rect 214 6071 662 6077
rect 214 6048 252 6071
rect 153 6034 252 6048
rect 153 5982 162 6034
rect 214 6019 252 6034
rect 304 6019 316 6071
rect 368 6019 380 6071
rect 432 6019 444 6071
rect 496 6019 508 6071
rect 560 6048 662 6071
rect 696 6068 776 6082
rect 696 6048 736 6068
rect 560 6034 736 6048
rect 770 6034 776 6068
rect 560 6019 776 6034
rect 214 6009 776 6019
rect 214 6002 662 6009
rect 214 5982 252 6002
rect 153 5968 252 5982
rect 153 5916 162 5968
rect 214 5950 252 5968
rect 304 5950 316 6002
rect 368 5950 380 6002
rect 432 5950 444 6002
rect 496 5950 508 6002
rect 560 5975 662 6002
rect 696 5996 776 6009
rect 696 5975 736 5996
rect 560 5962 736 5975
rect 770 5962 776 5996
rect 560 5950 776 5962
rect 214 5936 776 5950
rect 214 5933 662 5936
rect 214 5916 252 5933
rect 153 5902 252 5916
rect 153 5850 162 5902
rect 214 5881 252 5902
rect 304 5881 316 5933
rect 368 5881 380 5933
rect 432 5881 444 5933
rect 496 5881 508 5933
rect 560 5902 662 5933
rect 696 5924 776 5936
rect 696 5902 736 5924
rect 560 5890 736 5902
rect 770 5890 776 5924
rect 560 5881 776 5890
rect 214 5864 776 5881
rect 214 5850 252 5864
rect 153 5836 252 5850
rect 153 5784 162 5836
rect 214 5812 252 5836
rect 304 5812 316 5864
rect 368 5812 380 5864
rect 432 5812 444 5864
rect 496 5812 508 5864
rect 560 5863 776 5864
rect 560 5829 662 5863
rect 696 5852 776 5863
rect 696 5829 736 5852
rect 560 5818 736 5829
rect 770 5818 776 5852
rect 560 5812 776 5818
rect 214 5795 776 5812
rect 214 5784 252 5795
rect 153 5777 171 5784
rect 205 5777 252 5784
rect 153 5770 252 5777
rect 153 5718 162 5770
rect 214 5743 252 5770
rect 304 5743 316 5795
rect 368 5743 380 5795
rect 432 5743 444 5795
rect 496 5743 508 5795
rect 560 5790 776 5795
rect 560 5756 662 5790
rect 696 5780 776 5790
rect 696 5756 736 5780
rect 560 5746 736 5756
rect 770 5746 776 5780
rect 560 5743 776 5746
rect 214 5726 776 5743
rect 214 5718 252 5726
rect 153 5704 171 5718
rect 205 5704 252 5718
rect 153 5652 162 5704
rect 214 5674 252 5704
rect 304 5674 316 5726
rect 368 5674 380 5726
rect 432 5674 444 5726
rect 496 5674 508 5726
rect 560 5717 776 5726
rect 560 5683 662 5717
rect 696 5708 776 5717
rect 696 5683 736 5708
rect 560 5674 736 5683
rect 770 5674 776 5708
rect 214 5657 776 5674
rect 214 5652 252 5657
rect 153 5638 171 5652
rect 205 5638 252 5652
rect 153 5586 162 5638
rect 214 5605 252 5638
rect 304 5605 316 5657
rect 368 5605 380 5657
rect 432 5605 444 5657
rect 496 5605 508 5657
rect 560 5644 776 5657
rect 560 5610 662 5644
rect 696 5636 776 5644
rect 696 5610 736 5636
rect 560 5605 736 5610
rect 214 5602 736 5605
rect 770 5602 776 5636
rect 214 5588 776 5602
rect 214 5586 252 5588
rect 153 5572 171 5586
rect 205 5572 252 5586
rect 153 5520 162 5572
rect 214 5536 252 5572
rect 304 5536 316 5588
rect 368 5536 380 5588
rect 432 5536 444 5588
rect 496 5536 508 5588
rect 560 5571 776 5588
rect 560 5537 662 5571
rect 696 5564 776 5571
rect 696 5537 736 5564
rect 560 5536 736 5537
rect 214 5530 736 5536
rect 770 5530 776 5564
rect 214 5520 776 5530
rect 153 5519 776 5520
rect 153 5506 171 5519
rect 205 5506 252 5519
rect 153 5454 162 5506
rect 214 5467 252 5506
rect 304 5467 316 5519
rect 368 5467 380 5519
rect 432 5467 444 5519
rect 496 5467 508 5519
rect 560 5498 776 5519
rect 560 5467 662 5498
rect 214 5464 662 5467
rect 696 5492 776 5498
rect 696 5464 736 5492
rect 214 5458 736 5464
rect 770 5458 776 5492
rect 214 5454 776 5458
rect 153 5449 776 5454
rect 153 5446 252 5449
rect 153 5440 171 5446
rect 205 5440 252 5446
rect 153 5388 162 5440
rect 214 5397 252 5440
rect 304 5397 316 5449
rect 368 5397 380 5449
rect 432 5397 444 5449
rect 496 5397 508 5449
rect 560 5425 776 5449
rect 560 5397 662 5425
rect 214 5391 662 5397
rect 696 5420 776 5425
rect 696 5391 736 5420
rect 214 5388 736 5391
rect 153 5386 736 5388
rect 770 5386 776 5420
rect 153 5379 776 5386
rect 153 5374 252 5379
rect 153 5322 162 5374
rect 214 5327 252 5374
rect 304 5327 316 5379
rect 368 5327 380 5379
rect 432 5327 444 5379
rect 496 5327 508 5379
rect 560 5352 776 5379
rect 560 5327 662 5352
rect 214 5322 662 5327
rect 153 5318 662 5322
rect 696 5348 776 5352
rect 696 5318 736 5348
rect 153 5314 736 5318
rect 770 5314 776 5348
rect 153 5300 776 5314
rect 153 5266 171 5300
rect 205 5279 776 5300
rect 205 5266 662 5279
rect 153 5245 662 5266
rect 696 5275 776 5279
rect 696 5245 736 5275
rect 153 5241 736 5245
rect 770 5241 776 5275
rect 153 5227 776 5241
rect 153 5193 171 5227
rect 205 5207 776 5227
rect 205 5193 297 5207
rect 153 5173 297 5193
rect 331 5173 370 5207
rect 404 5173 443 5207
rect 477 5173 516 5207
rect 550 5173 589 5207
rect 623 5202 776 5207
rect 623 5173 736 5202
rect 153 5168 736 5173
rect 770 5168 776 5202
rect 153 5154 776 5168
rect 153 5120 171 5154
rect 205 5130 776 5154
rect 205 5120 297 5130
rect 153 5096 297 5120
rect 331 5096 371 5130
rect 405 5096 444 5130
rect 478 5096 517 5130
rect 551 5096 590 5130
rect 624 5096 663 5130
rect 697 5096 776 5130
rect 153 5090 776 5096
rect -26 5031 -20 5065
rect 14 5031 52 5065
rect 86 5031 92 5065
rect -26 5016 92 5031
rect -26 5010 952 5016
rect -26 4992 129 5010
rect -26 4958 -20 4992
rect 14 4958 52 4992
rect 86 4976 129 4992
rect 163 4976 205 5010
rect 239 4976 281 5010
rect 315 4976 357 5010
rect 391 4976 433 5010
rect 467 4976 508 5010
rect 542 4976 583 5010
rect 617 4976 658 5010
rect 692 4976 733 5010
rect 767 4976 808 5010
rect 842 4976 952 5010
rect 86 4970 952 4976
rect 86 4958 92 4970
rect -26 4919 92 4958
rect -26 4885 -20 4919
rect 14 4885 52 4919
rect 86 4885 92 4919
tri 824 4914 880 4970 ne
rect 880 4914 952 4970
rect -26 4846 92 4885
rect -26 4812 -20 4846
rect 14 4812 52 4846
rect 86 4812 92 4846
rect -26 4773 92 4812
rect -26 4739 -20 4773
rect 14 4739 52 4773
rect 86 4739 92 4773
rect -26 4700 92 4739
rect -26 4666 -20 4700
rect 14 4666 52 4700
rect 86 4666 92 4700
rect -26 4627 92 4666
rect -26 4593 -20 4627
rect 14 4593 52 4627
rect 86 4593 92 4627
rect -26 4554 92 4593
rect -26 4520 -20 4554
rect 14 4520 52 4554
rect 86 4520 92 4554
rect -26 4481 92 4520
rect -26 4447 -20 4481
rect 14 4447 52 4481
rect 86 4447 92 4481
rect -26 4408 92 4447
rect -26 4374 -20 4408
rect 14 4374 52 4408
rect 86 4374 92 4408
rect -26 4335 92 4374
rect -26 4301 -20 4335
rect 14 4301 52 4335
rect 86 4301 92 4335
rect -26 4262 92 4301
rect -26 4228 -20 4262
rect 14 4228 52 4262
rect 86 4228 92 4262
rect -26 4189 92 4228
rect -26 4155 -20 4189
rect 14 4155 52 4189
rect 86 4155 92 4189
rect -26 4116 92 4155
rect -26 4082 -20 4116
rect 14 4082 52 4116
rect 86 4082 92 4116
rect -26 4043 92 4082
rect -26 4009 -20 4043
rect 14 4009 52 4043
rect 86 4009 92 4043
rect -26 3970 92 4009
rect -26 3936 -20 3970
rect 14 3936 52 3970
rect 86 3936 92 3970
rect -26 3897 92 3936
rect -26 3863 -20 3897
rect 14 3863 52 3897
rect 86 3863 92 3897
rect -26 3824 92 3863
rect -26 3790 -20 3824
rect 14 3790 52 3824
rect 86 3790 92 3824
rect -26 3751 92 3790
rect -26 3717 -20 3751
rect 14 3717 52 3751
rect 86 3717 92 3751
rect -26 3678 92 3717
rect -26 3644 -20 3678
rect 14 3644 52 3678
rect 86 3644 92 3678
rect -26 3605 92 3644
rect -26 3571 -20 3605
rect 14 3571 52 3605
rect 86 3571 92 3605
rect -26 3532 92 3571
rect -26 3498 -20 3532
rect 14 3498 52 3532
rect 86 3498 92 3532
rect -26 3459 92 3498
rect -26 3425 -20 3459
rect 14 3425 52 3459
rect 86 3425 92 3459
rect -26 3386 92 3425
rect -26 3352 -20 3386
rect 14 3352 52 3386
rect 86 3352 92 3386
rect -26 3313 92 3352
rect -26 3279 -20 3313
rect 14 3279 52 3313
rect 86 3279 92 3313
rect -26 3240 92 3279
rect -26 3206 -20 3240
rect 14 3206 52 3240
rect 86 3206 92 3240
rect -26 3167 92 3206
rect -26 3133 -20 3167
rect 14 3133 52 3167
rect 86 3133 92 3167
tri -54 3097 -26 3125 se
rect -26 3097 92 3133
tri -57 3094 -54 3097 se
rect -54 3094 92 3097
tri -91 3060 -57 3094 se
rect -57 3060 -20 3094
rect 14 3060 52 3094
rect 86 3060 92 3094
tri -94 3057 -91 3060 se
rect -91 3057 92 3060
tri -128 3023 -94 3057 se
rect -94 3023 92 3057
tri -130 3021 -128 3023 se
rect -128 3021 92 3023
tri -164 2987 -130 3021 se
rect -130 2987 -20 3021
rect 14 2987 52 3021
rect 86 2987 92 3021
rect 153 4908 796 4914
rect 153 4906 272 4908
rect 153 4854 162 4906
rect 214 4874 272 4906
rect 306 4874 354 4908
rect 388 4874 436 4908
rect 470 4874 518 4908
rect 552 4874 601 4908
rect 635 4874 684 4908
rect 718 4874 796 4908
rect 214 4854 796 4874
tri 880 4870 924 4914 ne
rect 924 4870 952 4914
rect 153 4838 796 4854
rect 153 4786 162 4838
rect 214 4835 796 4838
rect 214 4820 756 4835
rect 214 4786 272 4820
rect 306 4786 351 4820
rect 385 4786 430 4820
rect 464 4786 509 4820
rect 543 4786 588 4820
rect 622 4786 668 4820
rect 702 4801 756 4820
rect 790 4801 796 4835
rect 702 4786 796 4801
rect 153 4770 796 4786
rect 153 4718 162 4770
rect 214 4762 796 4770
rect 214 4748 756 4762
rect 214 4718 668 4748
rect 153 4714 668 4718
rect 702 4728 756 4748
rect 790 4728 796 4762
rect 702 4714 796 4728
rect 153 4702 796 4714
rect 153 4650 162 4702
rect 214 4689 796 4702
rect 214 4676 756 4689
rect 214 4664 668 4676
rect 214 4650 252 4664
rect 304 4658 316 4664
rect 153 4647 171 4650
rect 205 4647 252 4650
rect 153 4634 252 4647
rect 153 4582 162 4634
rect 214 4612 252 4634
rect 304 4612 316 4624
rect 368 4612 380 4664
rect 432 4612 444 4664
rect 496 4612 508 4664
rect 560 4658 668 4664
rect 573 4642 668 4658
rect 702 4655 756 4676
rect 790 4655 796 4689
rect 702 4642 796 4655
rect 573 4624 796 4642
rect 560 4616 796 4624
rect 560 4612 756 4616
rect 214 4604 756 4612
rect 214 4590 668 4604
rect 214 4582 252 4590
rect 304 4583 316 4590
rect 153 4574 171 4582
rect 205 4574 252 4582
rect 153 4566 252 4574
rect 153 4514 162 4566
rect 214 4538 252 4566
rect 304 4538 316 4549
rect 368 4538 380 4590
rect 432 4538 444 4590
rect 496 4538 508 4590
rect 560 4583 668 4590
rect 573 4570 668 4583
rect 702 4582 756 4604
rect 790 4582 796 4616
rect 702 4570 796 4582
rect 573 4549 796 4570
rect 560 4543 796 4549
rect 560 4538 756 4543
rect 214 4532 756 4538
rect 214 4516 668 4532
rect 214 4514 252 4516
rect 153 4501 171 4514
rect 205 4501 252 4514
rect 304 4508 316 4516
rect 153 4498 252 4501
rect 153 4446 162 4498
rect 214 4464 252 4498
rect 304 4464 316 4474
rect 368 4464 380 4516
rect 432 4464 444 4516
rect 496 4464 508 4516
rect 560 4508 668 4516
rect 573 4498 668 4508
rect 702 4509 756 4532
rect 790 4509 796 4543
rect 702 4498 796 4509
rect 573 4474 796 4498
rect 560 4470 796 4474
rect 560 4464 756 4470
rect 214 4459 756 4464
rect 214 4446 668 4459
rect 153 4430 171 4446
rect 205 4442 668 4446
rect 205 4430 252 4442
rect 304 4433 316 4442
rect 153 4378 162 4430
rect 214 4390 252 4430
rect 304 4390 316 4399
rect 368 4390 380 4442
rect 432 4390 444 4442
rect 496 4390 508 4442
rect 560 4433 668 4442
rect 573 4425 668 4433
rect 702 4436 756 4459
rect 790 4436 796 4470
rect 702 4425 796 4436
rect 573 4399 796 4425
rect 560 4397 796 4399
rect 560 4390 756 4397
rect 214 4386 756 4390
rect 214 4378 668 4386
rect 153 4361 171 4378
rect 205 4368 668 4378
rect 205 4361 252 4368
rect 153 4309 162 4361
rect 214 4316 252 4361
rect 304 4357 316 4368
rect 304 4316 316 4323
rect 368 4316 380 4368
rect 432 4316 444 4368
rect 496 4316 508 4368
rect 560 4357 668 4368
rect 573 4352 668 4357
rect 702 4363 756 4386
rect 790 4363 796 4397
rect 702 4352 796 4363
rect 573 4324 796 4352
rect 573 4323 756 4324
rect 560 4316 756 4323
rect 214 4313 756 4316
rect 214 4309 668 4313
rect 153 4292 171 4309
rect 205 4294 668 4309
rect 205 4292 252 4294
rect 153 4240 162 4292
rect 214 4242 252 4292
rect 304 4281 316 4294
rect 304 4242 316 4247
rect 368 4242 380 4294
rect 432 4242 444 4294
rect 496 4242 508 4294
rect 560 4281 668 4294
rect 573 4279 668 4281
rect 702 4290 756 4313
rect 790 4290 796 4324
rect 702 4279 796 4290
rect 573 4251 796 4279
rect 573 4247 756 4251
rect 560 4242 756 4247
rect 214 4240 756 4242
rect 153 4223 171 4240
rect 205 4223 668 4240
rect 153 4171 162 4223
rect 214 4220 668 4223
rect 214 4171 252 4220
rect 304 4205 316 4220
rect 153 4168 252 4171
rect 304 4168 316 4171
rect 368 4168 380 4220
rect 432 4168 444 4220
rect 496 4168 508 4220
rect 560 4206 668 4220
rect 702 4217 756 4240
rect 790 4217 796 4251
rect 702 4206 796 4217
rect 560 4205 796 4206
rect 573 4178 796 4205
rect 573 4171 756 4178
rect 560 4168 756 4171
rect 153 4167 756 4168
rect 153 4133 171 4167
rect 205 4133 668 4167
rect 702 4144 756 4167
rect 790 4144 796 4178
rect 702 4133 796 4144
rect 153 4129 796 4133
rect 153 4095 284 4129
rect 318 4095 539 4129
rect 573 4105 796 4129
rect 573 4095 756 4105
rect 153 4094 756 4095
rect 153 4093 668 4094
rect 153 4059 171 4093
rect 205 4060 668 4093
rect 702 4071 756 4094
rect 790 4071 796 4105
rect 702 4060 796 4071
rect 205 4059 796 4060
rect 153 4053 796 4059
rect 153 4019 284 4053
rect 318 4019 539 4053
rect 573 4032 796 4053
rect 573 4021 756 4032
rect 573 4019 668 4021
rect 153 3985 171 4019
rect 205 3987 668 4019
rect 702 3998 756 4021
rect 790 3998 796 4032
rect 702 3987 796 3998
rect 205 3985 796 3987
rect 153 3977 796 3985
rect 153 3945 284 3977
rect 153 3911 171 3945
rect 205 3943 284 3945
rect 318 3943 539 3977
rect 573 3959 796 3977
rect 573 3948 756 3959
rect 573 3943 668 3948
rect 205 3914 668 3943
rect 702 3925 756 3948
rect 790 3925 796 3959
rect 702 3914 796 3925
rect 205 3911 796 3914
rect 153 3901 796 3911
rect 153 3871 284 3901
rect 153 3837 171 3871
rect 205 3867 284 3871
rect 318 3867 539 3901
rect 573 3886 796 3901
rect 573 3875 756 3886
rect 573 3867 668 3875
rect 205 3841 668 3867
rect 702 3852 756 3875
rect 790 3852 796 3886
rect 702 3841 796 3852
rect 205 3837 796 3841
rect 153 3825 796 3837
rect 153 3797 284 3825
rect 153 3763 171 3797
rect 205 3791 284 3797
rect 318 3791 539 3825
rect 573 3813 796 3825
rect 573 3802 756 3813
rect 573 3791 668 3802
rect 205 3779 668 3791
rect 205 3768 267 3779
tri 267 3768 278 3779 nw
rect 662 3768 668 3779
rect 702 3779 756 3802
rect 790 3779 796 3813
rect 702 3768 796 3779
rect 205 3763 239 3768
rect 153 3740 239 3763
tri 239 3740 267 3768 nw
rect 662 3740 796 3768
rect 153 3729 228 3740
tri 228 3729 239 3740 nw
rect 662 3729 756 3740
rect 153 3723 223 3729
tri 223 3724 228 3729 nw
rect 153 3689 171 3723
rect 205 3689 223 3723
rect 153 3649 223 3689
rect 153 3615 171 3649
rect 205 3615 223 3649
rect 153 3575 223 3615
rect 153 3541 171 3575
rect 205 3541 223 3575
rect 153 3501 223 3541
rect 153 3467 171 3501
rect 205 3467 223 3501
rect 662 3695 668 3729
rect 702 3706 756 3729
rect 790 3706 796 3740
rect 702 3695 796 3706
rect 662 3667 796 3695
rect 662 3656 756 3667
rect 662 3622 668 3656
rect 702 3633 756 3656
rect 790 3633 796 3667
rect 702 3622 796 3633
rect 662 3593 796 3622
rect 662 3583 756 3593
rect 662 3549 668 3583
rect 702 3559 756 3583
rect 790 3559 796 3593
rect 702 3549 796 3559
rect 662 3519 796 3549
rect 662 3510 756 3519
rect 153 3427 223 3467
rect 153 3393 171 3427
rect 205 3393 223 3427
rect 153 3353 223 3393
rect 153 3319 171 3353
rect 205 3319 223 3353
rect 153 3279 223 3319
rect 153 3276 171 3279
rect 205 3276 223 3279
rect 153 3224 162 3276
rect 214 3224 223 3276
rect 153 3207 223 3224
rect 153 3155 162 3207
rect 214 3155 223 3207
rect 153 3138 223 3155
rect 153 3086 162 3138
rect 214 3086 223 3138
rect 153 3069 223 3086
rect 153 3017 162 3069
rect 214 3017 223 3069
rect 153 3011 223 3017
rect 364 3467 410 3479
rect 364 3433 370 3467
rect 404 3433 410 3467
rect 364 3393 410 3433
rect 364 3359 370 3393
rect 404 3359 410 3393
rect 364 3319 410 3359
rect 364 3285 370 3319
rect 404 3285 410 3319
rect 364 3245 410 3285
rect 364 3211 370 3245
rect 404 3211 410 3245
rect 364 3171 410 3211
rect 364 3137 370 3171
rect 404 3137 410 3171
rect 364 3097 410 3137
rect 364 3063 370 3097
rect 404 3063 410 3097
rect 364 3023 410 3063
tri -166 2985 -164 2987 se
rect -164 2985 92 2987
rect -166 2975 92 2985
rect 364 2989 370 3023
rect 404 2989 410 3023
rect -166 2965 -81 2975
tri -81 2965 -71 2975 nw
rect -166 2950 -96 2965
tri -96 2950 -81 2965 nw
rect 364 2950 410 2989
rect -166 2741 -108 2950
tri -108 2938 -96 2950 nw
rect 364 2916 370 2950
rect 404 2916 410 2950
tri 343 2892 364 2913 se
rect 364 2892 410 2916
tri 339 2888 343 2892 se
rect 343 2888 410 2892
rect -50 2877 410 2888
rect -50 2843 370 2877
rect 404 2843 410 2877
rect -50 2804 410 2843
rect 662 3476 668 3510
rect 702 3485 756 3510
rect 790 3485 796 3519
rect 702 3476 796 3485
rect 662 3445 796 3476
rect 662 3437 756 3445
rect 662 3403 668 3437
rect 702 3411 756 3437
rect 790 3411 796 3445
rect 702 3403 796 3411
rect 662 3371 796 3403
rect 662 3364 756 3371
rect 662 3330 668 3364
rect 702 3337 756 3364
rect 790 3337 796 3371
rect 702 3330 796 3337
rect 662 3297 796 3330
rect 662 3291 756 3297
rect 662 3257 668 3291
rect 702 3263 756 3291
rect 790 3263 796 3297
rect 702 3257 796 3263
rect 662 3223 796 3257
rect 662 3218 756 3223
rect 662 3184 668 3218
rect 702 3189 756 3218
rect 790 3189 796 3223
rect 702 3184 796 3189
rect 662 3149 796 3184
rect 662 3145 756 3149
rect 662 3111 668 3145
rect 702 3115 756 3145
rect 790 3115 796 3149
rect 702 3111 796 3115
rect 662 3075 796 3111
rect 662 3072 756 3075
rect 662 3038 668 3072
rect 702 3041 756 3072
rect 790 3041 796 3075
rect 702 3038 796 3041
rect 662 3001 796 3038
rect 662 2999 756 3001
rect 662 2965 668 2999
rect 702 2967 756 2999
rect 790 2967 796 3001
rect 702 2965 796 2967
rect 662 2927 796 2965
rect 662 2926 756 2927
rect 662 2892 668 2926
rect 702 2893 756 2926
rect 790 2893 796 2927
rect 702 2892 796 2893
rect 662 2853 796 2892
rect 662 2819 668 2853
rect 702 2819 756 2853
rect 790 2819 796 2853
rect 662 2807 796 2819
rect -50 2770 370 2804
rect 404 2770 410 2804
rect -50 2758 410 2770
rect 750 2775 796 2807
tri -108 2741 -105 2744 sw
rect 750 2741 756 2775
rect 790 2741 796 2775
rect -166 2716 -105 2741
tri -105 2716 -80 2741 sw
rect -166 2704 64 2716
rect -166 2670 -3 2704
rect 31 2670 64 2704
rect -166 2632 64 2670
tri -166 2598 -132 2632 ne
rect -132 2598 -3 2632
rect 31 2598 64 2632
tri -132 2593 -127 2598 ne
rect -127 2593 64 2598
tri -127 2587 -121 2593 ne
rect -121 2587 64 2593
tri -121 2560 -94 2587 ne
rect -94 2560 64 2587
tri -94 2526 -60 2560 ne
rect -60 2526 -3 2560
rect 31 2526 64 2560
tri -60 2517 -51 2526 ne
rect -51 2517 64 2526
tri -51 2510 -44 2517 ne
rect -44 2510 64 2517
tri -44 2505 -39 2510 ne
rect -39 2505 64 2510
rect 158 2702 306 2714
rect 158 2668 164 2702
rect 158 2650 167 2668
rect 219 2650 245 2702
rect 300 2668 306 2702
rect 297 2650 306 2668
rect 158 2635 306 2650
rect 158 2627 167 2635
rect 158 2593 164 2627
rect 158 2583 167 2593
rect 219 2583 245 2635
rect 297 2627 306 2635
rect 300 2593 306 2627
rect 297 2583 306 2593
rect 158 2568 306 2583
rect 158 2551 167 2568
rect 158 2517 164 2551
rect 158 2516 167 2517
rect 219 2516 245 2568
rect 297 2551 306 2568
rect 300 2517 306 2551
rect 297 2516 306 2517
rect 158 2505 306 2516
rect 750 2698 796 2741
rect 750 2664 756 2698
rect 790 2664 796 2698
rect 750 2621 796 2664
rect 750 2587 756 2621
rect 790 2587 796 2621
rect 750 2544 796 2587
rect 750 2510 756 2544
rect 790 2510 796 2544
tri -39 2502 -36 2505 ne
rect -36 2488 64 2505
rect -36 2454 -3 2488
rect 31 2454 64 2488
rect 750 2467 796 2510
rect -36 2416 64 2454
rect -36 2382 -3 2416
rect 31 2382 64 2416
rect -36 2344 64 2382
rect -36 2310 -3 2344
rect 31 2310 64 2344
rect 124 2446 512 2458
rect 124 2412 472 2446
rect 506 2412 512 2446
rect 124 2374 512 2412
rect 124 2340 472 2374
rect 506 2340 512 2374
rect 124 2328 512 2340
rect 750 2433 756 2467
rect 790 2433 796 2467
rect 750 2390 796 2433
rect 750 2356 756 2390
rect 790 2356 796 2390
rect -36 2271 64 2310
rect 750 2313 796 2356
rect -36 2237 -3 2271
rect 31 2237 64 2271
tri -53 2202 -36 2219 se
rect -36 2202 64 2237
tri -57 2198 -53 2202 se
rect -53 2198 64 2202
tri -91 2164 -57 2198 se
rect -57 2164 -3 2198
rect 31 2164 64 2198
tri -94 2161 -91 2164 se
rect -91 2161 64 2164
tri -97 2158 -94 2161 se
rect -94 2158 64 2161
tri -130 2125 -97 2158 se
rect -97 2125 64 2158
tri -164 2091 -130 2125 se
rect -130 2091 -3 2125
rect 31 2091 64 2125
tri -166 2089 -164 2091 se
rect -164 2089 64 2091
rect -166 2079 64 2089
rect 158 2270 306 2282
rect 158 2236 164 2270
rect 158 2218 167 2236
rect 219 2218 245 2270
rect 300 2236 306 2270
rect 297 2218 306 2236
rect 158 2203 306 2218
rect 158 2195 167 2203
rect 158 2161 164 2195
rect 158 2151 167 2161
rect 219 2151 245 2203
rect 297 2195 306 2203
rect 300 2161 306 2195
rect 297 2151 306 2161
rect 158 2136 306 2151
rect 158 2119 167 2136
rect 158 2085 164 2119
rect 158 2084 167 2085
rect 219 2084 245 2136
rect 297 2119 306 2136
rect 300 2085 306 2119
rect 297 2084 306 2085
rect -166 2073 -77 2079
tri -77 2073 -71 2079 nw
rect 158 2073 306 2084
rect 750 2279 756 2313
rect 790 2279 796 2313
rect 750 2236 796 2279
rect 750 2202 756 2236
rect 790 2202 796 2236
rect 750 2158 796 2202
rect 750 2124 756 2158
rect 790 2124 796 2158
rect 750 2080 796 2124
rect -166 2046 -104 2073
tri -104 2046 -77 2073 nw
rect 750 2046 756 2080
rect 790 2046 796 2080
rect -166 1834 -108 2046
tri -108 2042 -104 2046 nw
rect -50 2016 410 2028
rect -50 1982 370 2016
rect 404 1982 410 2016
rect -50 1942 410 1982
rect -50 1908 370 1942
rect 404 1908 410 1942
rect 750 2002 796 2046
rect 750 1968 756 2002
rect 790 1968 796 2002
rect 750 1936 796 1968
rect -50 1898 410 1908
tri 339 1890 347 1898 ne
rect 347 1890 410 1898
tri 347 1873 364 1890 ne
rect 364 1868 410 1890
tri -108 1834 -94 1848 sw
rect 364 1834 370 1868
rect 404 1834 410 1868
rect -166 1820 -94 1834
tri -94 1820 -80 1834 sw
rect -166 1808 68 1820
rect -166 1774 -44 1808
rect -10 1774 28 1808
rect 62 1774 68 1808
rect 364 1794 410 1834
rect -166 1736 68 1774
tri -166 1735 -165 1736 ne
rect -165 1735 28 1736
tri -165 1701 -131 1735 ne
rect -131 1701 -44 1735
rect -10 1702 28 1735
rect 62 1702 68 1736
rect -10 1701 68 1702
tri -131 1691 -121 1701 ne
rect -121 1691 68 1701
tri -121 1690 -120 1691 ne
rect -120 1690 68 1691
tri -120 1664 -94 1690 ne
rect -94 1664 68 1690
tri -94 1662 -92 1664 ne
rect -92 1662 28 1664
tri -92 1628 -58 1662 ne
rect -58 1628 -44 1662
rect -10 1630 28 1662
rect 62 1630 68 1664
rect -10 1628 68 1630
tri -58 1620 -50 1628 ne
rect -50 1592 68 1628
rect -50 1589 28 1592
rect -50 1555 -44 1589
rect -10 1558 28 1589
rect 62 1558 68 1592
rect -10 1555 68 1558
rect -50 1520 68 1555
rect -50 1516 28 1520
rect -50 1482 -44 1516
rect -10 1486 28 1516
rect 62 1486 68 1520
rect -10 1482 68 1486
rect -50 1448 68 1482
rect -50 1443 28 1448
rect -50 1409 -44 1443
rect -10 1414 28 1443
rect 62 1414 68 1448
rect 161 1764 295 1776
rect 161 1730 167 1764
rect 201 1730 255 1764
rect 289 1730 295 1764
rect 161 1691 295 1730
rect 161 1690 255 1691
rect 161 1656 167 1690
rect 201 1657 255 1690
rect 289 1657 295 1691
rect 201 1656 295 1657
rect 161 1618 295 1656
rect 161 1616 255 1618
rect 161 1582 167 1616
rect 201 1584 255 1616
rect 289 1584 295 1618
rect 201 1582 295 1584
rect 161 1545 295 1582
rect 161 1542 255 1545
rect 161 1508 167 1542
rect 201 1511 255 1542
rect 289 1511 295 1545
rect 201 1508 295 1511
rect 161 1472 295 1508
rect 161 1468 255 1472
rect 161 1434 167 1468
rect 201 1438 255 1468
rect 289 1438 295 1472
rect 201 1434 295 1438
rect 161 1424 295 1434
rect 364 1760 370 1794
rect 404 1760 410 1794
rect 364 1720 410 1760
rect 364 1686 370 1720
rect 404 1686 410 1720
rect 364 1646 410 1686
rect 364 1612 370 1646
rect 404 1612 410 1646
rect 364 1572 410 1612
rect 364 1538 370 1572
rect 404 1538 410 1572
rect 364 1498 410 1538
rect 364 1464 370 1498
rect 404 1464 410 1498
tri 295 1424 301 1430 sw
rect 364 1424 410 1464
rect -10 1409 68 1414
rect -50 1376 68 1409
rect -50 1370 28 1376
rect -50 1336 -44 1370
rect -10 1342 28 1370
rect 62 1342 68 1376
rect -10 1336 68 1342
rect -50 1304 68 1336
rect -50 1297 28 1304
rect -50 1263 -44 1297
rect -10 1270 28 1297
rect 62 1270 68 1304
rect -10 1263 68 1270
rect -50 1232 68 1263
rect -50 1224 28 1232
rect -50 1190 -44 1224
rect -10 1198 28 1224
rect 62 1198 68 1232
rect -10 1190 68 1198
rect -50 1160 68 1190
rect -50 1151 28 1160
rect -50 1117 -44 1151
rect -10 1126 28 1151
rect 62 1126 68 1160
rect -10 1117 68 1126
rect -50 1088 68 1117
rect -50 1077 28 1088
rect -50 1043 -44 1077
rect -10 1054 28 1077
rect 62 1054 68 1088
rect -10 1043 68 1054
rect -50 1016 68 1043
rect -50 1003 28 1016
rect -50 969 -44 1003
rect -10 982 28 1003
rect 62 982 68 1016
rect -10 969 68 982
rect -50 944 68 969
rect -50 929 28 944
rect -50 895 -44 929
rect -10 910 28 929
rect 62 910 68 944
rect -10 895 68 910
rect -50 872 68 895
rect -50 855 28 872
rect -50 821 -44 855
rect -10 838 28 855
rect 62 838 68 872
rect -10 821 68 838
tri 160 1415 161 1416 se
rect 161 1415 301 1424
tri 301 1415 310 1424 sw
rect 160 1409 310 1415
rect 212 1399 258 1409
rect 212 1365 255 1399
rect 212 1357 258 1365
rect 160 1344 310 1357
rect 212 1326 258 1344
rect 212 1292 255 1326
rect 160 1286 167 1292
rect 201 1286 310 1292
rect 160 1279 310 1286
rect 212 1253 258 1279
rect 212 1227 255 1253
rect 160 1214 167 1227
rect 201 1219 255 1227
rect 289 1219 310 1227
rect 201 1214 310 1219
rect 212 1180 258 1214
rect 212 1162 255 1180
rect 160 1149 167 1162
rect 201 1149 255 1162
rect 289 1149 310 1162
rect 212 1146 255 1149
rect 212 1107 258 1146
rect 212 1097 255 1107
rect 160 1084 167 1097
rect 201 1084 255 1097
rect 289 1084 310 1097
rect 212 1073 255 1084
rect 212 1034 258 1073
rect 212 1032 255 1034
rect 160 1025 255 1032
rect 160 1018 167 1025
rect 201 1018 255 1025
rect 289 1018 310 1032
rect 212 1000 255 1018
rect 212 966 258 1000
rect 160 961 310 966
rect 160 952 255 961
rect 289 952 310 961
rect 212 927 255 952
rect 212 900 258 927
rect 160 888 310 900
rect 160 886 255 888
rect 289 886 310 888
rect 212 854 255 886
rect 212 834 258 854
rect 160 828 310 834
tri 160 827 161 828 ne
rect -50 800 68 821
rect -50 781 28 800
rect -50 747 -44 781
rect -10 766 28 781
rect 62 766 68 800
rect -10 747 68 766
rect -50 728 68 747
rect -50 707 28 728
rect -50 673 -44 707
rect -10 694 28 707
rect 62 694 68 728
rect -10 673 68 694
rect -50 656 68 673
rect -50 633 28 656
rect -50 599 -44 633
rect -10 622 28 633
rect 62 622 68 656
rect -10 599 68 622
rect -50 584 68 599
rect -50 559 28 584
rect -50 525 -44 559
rect -10 550 28 559
rect 62 550 68 584
rect -10 525 68 550
rect -50 512 68 525
rect -50 485 28 512
rect -50 451 -44 485
rect -10 478 28 485
rect 62 478 68 512
rect -10 451 68 478
rect -50 440 68 451
rect -50 411 28 440
rect -50 377 -44 411
rect -10 406 28 411
rect 62 406 68 440
rect -10 377 68 406
rect -50 368 68 377
rect -50 337 28 368
rect -50 303 -44 337
rect -10 334 28 337
rect 62 334 68 368
rect -10 303 68 334
rect -50 296 68 303
rect -50 263 28 296
rect -50 229 -44 263
rect -10 262 28 263
rect 62 262 68 296
rect -10 229 68 262
rect -50 223 68 229
rect -50 189 28 223
rect 62 189 68 223
rect -50 155 -44 189
rect -10 155 68 189
rect 161 815 295 828
rect 161 806 255 815
rect 161 772 167 806
rect 201 781 255 806
rect 289 781 295 815
tri 295 813 310 828 nw
rect 364 1390 370 1424
rect 404 1390 410 1424
rect 364 1350 410 1390
rect 364 1316 370 1350
rect 404 1316 410 1350
rect 364 1276 410 1316
rect 364 1242 370 1276
rect 404 1242 410 1276
rect 364 1202 410 1242
rect 364 1168 370 1202
rect 404 1168 410 1202
rect 364 1129 410 1168
rect 364 1095 370 1129
rect 404 1095 410 1129
rect 364 1056 410 1095
rect 364 1022 370 1056
rect 404 1022 410 1056
rect 364 983 410 1022
rect 364 949 370 983
rect 404 949 410 983
rect 364 910 410 949
rect 364 876 370 910
rect 404 876 410 910
rect 364 837 410 876
rect 201 772 295 781
rect 161 742 295 772
rect 161 733 255 742
rect 161 699 167 733
rect 201 708 255 733
rect 289 708 295 742
rect 364 803 370 837
rect 404 803 410 837
rect 364 764 410 803
rect 364 730 370 764
rect 404 730 410 764
rect 364 718 410 730
rect 662 1924 796 1936
rect 662 1890 668 1924
rect 702 1890 756 1924
rect 790 1890 796 1924
rect 662 1851 796 1890
rect 662 1817 668 1851
rect 702 1850 796 1851
rect 702 1817 756 1850
rect 662 1816 756 1817
rect 790 1816 796 1850
rect 662 1778 796 1816
rect 662 1744 668 1778
rect 702 1776 796 1778
rect 702 1744 756 1776
rect 662 1742 756 1744
rect 790 1742 796 1776
rect 662 1705 796 1742
rect 662 1671 668 1705
rect 702 1702 796 1705
rect 702 1671 756 1702
rect 662 1668 756 1671
rect 790 1668 796 1702
rect 662 1632 796 1668
rect 662 1598 668 1632
rect 702 1628 796 1632
rect 702 1598 756 1628
rect 662 1594 756 1598
rect 790 1594 796 1628
rect 662 1559 796 1594
rect 662 1525 668 1559
rect 702 1554 796 1559
rect 702 1525 756 1554
rect 662 1520 756 1525
rect 790 1520 796 1554
rect 662 1486 796 1520
rect 662 1452 668 1486
rect 702 1480 796 1486
rect 702 1452 756 1480
rect 662 1446 756 1452
rect 790 1446 796 1480
rect 662 1413 796 1446
rect 662 1379 668 1413
rect 702 1406 796 1413
rect 702 1379 756 1406
rect 662 1372 756 1379
rect 790 1372 796 1406
rect 662 1340 796 1372
rect 662 1306 668 1340
rect 702 1332 796 1340
rect 702 1306 756 1332
rect 662 1298 756 1306
rect 790 1298 796 1332
rect 662 1267 796 1298
rect 662 1233 668 1267
rect 702 1258 796 1267
rect 702 1233 756 1258
rect 662 1224 756 1233
rect 790 1224 796 1258
rect 662 1194 796 1224
rect 662 1160 668 1194
rect 702 1184 796 1194
rect 702 1160 756 1184
rect 662 1150 756 1160
rect 790 1150 796 1184
rect 662 1121 796 1150
rect 662 1087 668 1121
rect 702 1110 796 1121
rect 702 1087 756 1110
rect 662 1076 756 1087
rect 790 1076 796 1110
rect 662 1048 796 1076
rect 662 1014 668 1048
rect 702 1036 796 1048
rect 702 1014 756 1036
rect 662 1002 756 1014
rect 790 1002 796 1036
rect 662 975 796 1002
rect 662 941 668 975
rect 702 962 796 975
rect 702 941 756 962
rect 662 928 756 941
rect 790 928 796 962
rect 662 902 796 928
rect 662 868 668 902
rect 702 888 796 902
rect 702 868 756 888
rect 662 854 756 868
rect 790 854 796 888
rect 662 828 796 854
rect 662 794 668 828
rect 702 814 796 828
rect 702 794 756 814
rect 662 780 756 794
rect 790 780 796 814
rect 662 754 796 780
rect 662 720 668 754
rect 702 740 796 754
rect 702 720 756 740
rect 201 699 295 708
rect 161 670 295 699
rect 161 660 255 670
rect 161 626 167 660
rect 201 636 255 660
rect 289 636 295 670
rect 201 626 295 636
rect 161 598 295 626
rect 161 587 255 598
rect 161 553 167 587
rect 201 564 255 587
rect 289 564 295 598
rect 201 553 295 564
rect 161 526 295 553
rect 161 514 255 526
rect 161 480 167 514
rect 201 492 255 514
rect 289 492 295 526
rect 201 480 295 492
rect 161 454 295 480
rect 161 441 255 454
rect 161 407 167 441
rect 201 420 255 441
rect 289 420 295 454
rect 662 706 756 720
rect 790 706 796 740
rect 662 680 796 706
rect 662 646 668 680
rect 702 666 796 680
rect 702 646 756 666
rect 662 632 756 646
rect 790 632 796 666
rect 662 606 796 632
rect 662 572 668 606
rect 702 592 796 606
rect 702 572 756 592
rect 662 558 756 572
rect 790 558 796 592
rect 662 532 796 558
rect 662 498 668 532
rect 702 518 796 532
rect 702 498 756 518
rect 662 484 756 498
rect 790 484 796 518
rect 662 458 796 484
rect 662 424 668 458
rect 702 444 796 458
rect 702 424 756 444
rect 201 410 295 420
tri 295 410 308 423 sw
tri 649 410 662 423 se
rect 662 410 756 424
rect 790 410 796 444
rect 201 407 308 410
rect 161 384 308 407
tri 308 384 334 410 sw
tri 623 384 649 410 se
rect 649 384 796 410
rect 161 382 334 384
rect 161 368 255 382
rect 161 334 167 368
rect 201 348 255 368
rect 289 350 334 382
tri 334 350 368 384 sw
tri 589 350 623 384 se
rect 623 350 668 384
rect 702 369 796 384
rect 702 350 756 369
rect 289 348 368 350
rect 201 335 368 348
tri 368 335 383 350 sw
tri 574 335 589 350 se
rect 589 335 756 350
rect 790 335 796 369
rect 201 334 383 335
rect 161 316 383 334
tri 383 316 402 335 sw
tri 555 316 574 335 se
rect 574 316 796 335
rect 161 310 796 316
rect 161 295 255 310
rect 161 261 167 295
rect 201 276 255 295
rect 289 276 338 310
rect 372 276 421 310
rect 455 276 504 310
rect 538 276 586 310
rect 620 276 668 310
rect 702 294 796 310
rect 702 276 756 294
rect 201 261 756 276
rect 161 260 756 261
rect 790 260 796 294
rect 161 222 796 260
rect 161 188 239 222
rect 273 188 313 222
rect 347 188 387 222
rect 421 188 461 222
rect 495 188 535 222
rect 569 188 609 222
rect 643 188 683 222
rect 717 188 796 222
rect 161 182 796 188
tri 857 182 908 233 se
rect 908 182 1149 233
tri 852 177 857 182 se
rect 857 177 1149 182
rect -50 115 68 155
rect -50 81 -44 115
rect -10 107 68 115
tri 68 107 138 177 sw
tri 782 107 852 177 se
rect 852 167 1149 177
rect 852 107 1089 167
tri 1089 107 1149 167 nw
rect -10 101 1043 107
rect -10 81 59 101
rect -50 67 59 81
rect 93 67 134 101
rect 168 67 209 101
rect 243 67 284 101
rect 318 67 359 101
rect 393 67 434 101
rect 468 67 509 101
rect 543 67 584 101
rect 618 67 659 101
rect 693 67 734 101
rect 768 67 808 101
rect 842 67 1043 101
rect -50 61 1043 67
tri 1043 61 1089 107 nw
rect -50 41 936 61
rect -50 7 -44 41
rect -10 7 936 41
rect -50 -46 936 7
tri 936 -46 1043 61 nw
<< via1 >>
rect 154 10281 206 10292
rect 154 10247 158 10281
rect 158 10247 192 10281
rect 192 10247 206 10281
rect 154 10240 206 10247
rect 258 10281 310 10292
rect 258 10247 278 10281
rect 278 10247 310 10281
rect 258 10240 310 10247
rect 154 10168 158 10188
rect 158 10168 192 10188
rect 192 10168 206 10188
rect 154 10136 206 10168
rect 258 10168 278 10188
rect 278 10168 310 10188
rect 258 10136 310 10168
rect 154 10043 206 10083
rect 154 10031 158 10043
rect 158 10031 192 10043
rect 192 10031 206 10043
rect 258 10043 310 10083
rect 258 10031 278 10043
rect 278 10031 310 10043
rect 154 9963 206 9978
rect 154 9929 158 9963
rect 158 9929 192 9963
rect 192 9929 206 9963
rect 154 9926 206 9929
rect 258 9963 310 9978
rect 258 9929 278 9963
rect 278 9929 310 9963
rect 258 9926 310 9929
rect 154 9849 158 9873
rect 158 9849 192 9873
rect 192 9849 206 9873
rect 154 9821 206 9849
rect 258 9849 278 9873
rect 278 9849 310 9873
rect 258 9821 310 9849
rect 154 9716 206 9768
rect 258 9716 310 9768
rect 154 8463 206 8477
rect 154 8429 158 8463
rect 158 8429 192 8463
rect 192 8429 206 8463
rect 154 8425 206 8429
rect 258 8463 310 8477
rect 258 8429 278 8463
rect 278 8429 310 8463
rect 258 8425 310 8429
rect 154 8384 206 8412
rect 154 8360 158 8384
rect 158 8360 192 8384
rect 192 8360 206 8384
rect 258 8384 310 8412
rect 258 8360 278 8384
rect 278 8360 310 8384
rect 154 8305 206 8347
rect 154 8295 158 8305
rect 158 8295 192 8305
rect 192 8295 206 8305
rect 258 8305 310 8347
rect 258 8295 278 8305
rect 278 8295 310 8305
rect 154 8271 158 8282
rect 158 8271 192 8282
rect 192 8271 206 8282
rect 154 8230 206 8271
rect 258 8271 278 8282
rect 278 8271 310 8282
rect 258 8230 310 8271
rect 154 8191 158 8217
rect 158 8191 192 8217
rect 192 8191 206 8217
rect 154 8165 206 8191
rect 258 8191 278 8217
rect 278 8191 310 8217
rect 258 8165 310 8191
rect 154 8145 206 8151
rect 154 8111 158 8145
rect 158 8111 192 8145
rect 192 8111 206 8145
rect 154 8099 206 8111
rect 258 8145 310 8151
rect 258 8111 278 8145
rect 278 8111 310 8145
rect 258 8099 310 8111
rect 154 8065 206 8085
rect 154 8033 158 8065
rect 158 8033 192 8065
rect 192 8033 206 8065
rect 258 8065 310 8085
rect 258 8033 278 8065
rect 278 8033 310 8065
rect 154 7967 206 8019
rect 258 7967 310 8019
rect 154 7901 206 7953
rect 258 7901 310 7953
rect 162 7052 214 7087
rect 162 7035 171 7052
rect 171 7035 205 7052
rect 205 7035 214 7052
rect 162 7018 171 7022
rect 171 7018 205 7022
rect 205 7018 214 7022
rect 162 6979 214 7018
rect 162 6970 171 6979
rect 171 6970 205 6979
rect 205 6970 214 6979
rect 162 6945 171 6957
rect 171 6945 205 6957
rect 205 6945 214 6957
rect 162 6906 214 6945
rect 162 6905 171 6906
rect 171 6905 205 6906
rect 205 6905 214 6906
rect 162 6872 171 6892
rect 171 6872 205 6892
rect 205 6872 214 6892
rect 162 6840 214 6872
rect 162 6799 171 6826
rect 171 6799 205 6826
rect 205 6799 214 6826
rect 162 6774 214 6799
rect 162 6726 171 6760
rect 171 6726 205 6760
rect 205 6726 214 6760
rect 162 6708 214 6726
rect 162 6687 214 6694
rect 162 6653 171 6687
rect 171 6653 205 6687
rect 205 6653 214 6687
rect 162 6642 214 6653
rect 162 6614 214 6628
rect 162 6580 171 6614
rect 171 6580 205 6614
rect 205 6580 214 6614
rect 162 6576 214 6580
rect 162 6541 214 6562
rect 162 6510 171 6541
rect 171 6510 205 6541
rect 205 6510 214 6541
rect 162 6468 214 6496
rect 162 6444 171 6468
rect 171 6444 205 6468
rect 205 6444 214 6468
rect 162 6395 214 6430
rect 162 6378 171 6395
rect 171 6378 205 6395
rect 205 6378 214 6395
rect 162 6361 171 6364
rect 171 6361 205 6364
rect 205 6361 214 6364
rect 162 6322 214 6361
rect 162 6312 171 6322
rect 171 6312 205 6322
rect 205 6312 214 6322
rect 162 6288 171 6298
rect 171 6288 205 6298
rect 205 6288 214 6298
rect 162 6249 214 6288
rect 162 6246 171 6249
rect 171 6246 205 6249
rect 205 6246 214 6249
rect 162 6215 171 6232
rect 171 6215 205 6232
rect 205 6215 214 6232
rect 162 6180 214 6215
rect 162 6142 171 6166
rect 171 6142 205 6166
rect 205 6142 214 6166
rect 162 6114 214 6142
rect 162 6069 171 6100
rect 171 6069 205 6100
rect 205 6069 214 6100
rect 162 6048 214 6069
rect 162 6030 214 6034
rect 162 5996 171 6030
rect 171 5996 205 6030
rect 205 5996 214 6030
rect 252 6019 304 6071
rect 316 6019 368 6071
rect 380 6019 432 6071
rect 444 6019 496 6071
rect 508 6019 560 6071
rect 162 5982 214 5996
rect 162 5957 214 5968
rect 162 5923 171 5957
rect 171 5923 205 5957
rect 205 5923 214 5957
rect 252 5950 304 6002
rect 316 5950 368 6002
rect 380 5950 432 6002
rect 444 5950 496 6002
rect 508 5950 560 6002
rect 162 5916 214 5923
rect 162 5884 214 5902
rect 162 5850 171 5884
rect 171 5850 205 5884
rect 205 5850 214 5884
rect 252 5881 304 5933
rect 316 5881 368 5933
rect 380 5881 432 5933
rect 444 5881 496 5933
rect 508 5881 560 5933
rect 162 5811 214 5836
rect 252 5812 304 5864
rect 316 5812 368 5864
rect 380 5812 432 5864
rect 444 5812 496 5864
rect 508 5812 560 5864
rect 162 5784 171 5811
rect 171 5784 205 5811
rect 205 5784 214 5811
rect 162 5738 214 5770
rect 252 5743 304 5795
rect 316 5743 368 5795
rect 380 5743 432 5795
rect 444 5743 496 5795
rect 508 5743 560 5795
rect 162 5718 171 5738
rect 171 5718 205 5738
rect 205 5718 214 5738
rect 162 5665 214 5704
rect 252 5674 304 5726
rect 316 5674 368 5726
rect 380 5674 432 5726
rect 444 5674 496 5726
rect 508 5674 560 5726
rect 162 5652 171 5665
rect 171 5652 205 5665
rect 205 5652 214 5665
rect 162 5631 171 5638
rect 171 5631 205 5638
rect 205 5631 214 5638
rect 162 5592 214 5631
rect 252 5605 304 5657
rect 316 5605 368 5657
rect 380 5605 432 5657
rect 444 5605 496 5657
rect 508 5605 560 5657
rect 162 5586 171 5592
rect 171 5586 205 5592
rect 205 5586 214 5592
rect 162 5558 171 5572
rect 171 5558 205 5572
rect 205 5558 214 5572
rect 162 5520 214 5558
rect 252 5536 304 5588
rect 316 5536 368 5588
rect 380 5536 432 5588
rect 444 5536 496 5588
rect 508 5536 560 5588
rect 162 5485 171 5506
rect 171 5485 205 5506
rect 205 5485 214 5506
rect 162 5454 214 5485
rect 252 5467 304 5519
rect 316 5467 368 5519
rect 380 5467 432 5519
rect 444 5467 496 5519
rect 508 5467 560 5519
rect 162 5412 171 5440
rect 171 5412 205 5440
rect 205 5412 214 5440
rect 162 5388 214 5412
rect 252 5397 304 5449
rect 316 5397 368 5449
rect 380 5397 432 5449
rect 444 5397 496 5449
rect 508 5397 560 5449
rect 162 5373 214 5374
rect 162 5339 171 5373
rect 171 5339 205 5373
rect 205 5339 214 5373
rect 162 5322 214 5339
rect 252 5327 304 5379
rect 316 5327 368 5379
rect 380 5327 432 5379
rect 444 5327 496 5379
rect 508 5327 560 5379
rect 162 4900 214 4906
rect 162 4866 171 4900
rect 171 4866 205 4900
rect 205 4866 214 4900
rect 162 4854 214 4866
rect 162 4827 214 4838
rect 162 4793 171 4827
rect 171 4793 205 4827
rect 205 4793 214 4827
rect 162 4786 214 4793
rect 162 4754 214 4770
rect 162 4720 171 4754
rect 171 4720 205 4754
rect 205 4720 214 4754
rect 162 4718 214 4720
rect 162 4681 214 4702
rect 162 4650 171 4681
rect 171 4650 205 4681
rect 205 4650 214 4681
rect 252 4658 304 4664
rect 316 4658 368 4664
rect 162 4608 214 4634
rect 252 4624 284 4658
rect 284 4624 304 4658
rect 316 4624 318 4658
rect 318 4624 368 4658
rect 252 4612 304 4624
rect 316 4612 368 4624
rect 380 4612 432 4664
rect 444 4612 496 4664
rect 508 4658 560 4664
rect 508 4624 539 4658
rect 539 4624 560 4658
rect 508 4612 560 4624
rect 162 4582 171 4608
rect 171 4582 205 4608
rect 205 4582 214 4608
rect 252 4583 304 4590
rect 316 4583 368 4590
rect 162 4535 214 4566
rect 252 4549 284 4583
rect 284 4549 304 4583
rect 316 4549 318 4583
rect 318 4549 368 4583
rect 252 4538 304 4549
rect 316 4538 368 4549
rect 380 4538 432 4590
rect 444 4538 496 4590
rect 508 4583 560 4590
rect 508 4549 539 4583
rect 539 4549 560 4583
rect 508 4538 560 4549
rect 162 4514 171 4535
rect 171 4514 205 4535
rect 205 4514 214 4535
rect 252 4508 304 4516
rect 316 4508 368 4516
rect 162 4462 214 4498
rect 252 4474 284 4508
rect 284 4474 304 4508
rect 316 4474 318 4508
rect 318 4474 368 4508
rect 252 4464 304 4474
rect 316 4464 368 4474
rect 380 4464 432 4516
rect 444 4464 496 4516
rect 508 4508 560 4516
rect 508 4474 539 4508
rect 539 4474 560 4508
rect 508 4464 560 4474
rect 162 4446 171 4462
rect 171 4446 205 4462
rect 205 4446 214 4462
rect 252 4433 304 4442
rect 316 4433 368 4442
rect 162 4428 171 4430
rect 171 4428 205 4430
rect 205 4428 214 4430
rect 162 4389 214 4428
rect 252 4399 284 4433
rect 284 4399 304 4433
rect 316 4399 318 4433
rect 318 4399 368 4433
rect 252 4390 304 4399
rect 316 4390 368 4399
rect 380 4390 432 4442
rect 444 4390 496 4442
rect 508 4433 560 4442
rect 508 4399 539 4433
rect 539 4399 560 4433
rect 508 4390 560 4399
rect 162 4378 171 4389
rect 171 4378 205 4389
rect 205 4378 214 4389
rect 162 4355 171 4361
rect 171 4355 205 4361
rect 205 4355 214 4361
rect 162 4315 214 4355
rect 252 4357 304 4368
rect 316 4357 368 4368
rect 252 4323 284 4357
rect 284 4323 304 4357
rect 316 4323 318 4357
rect 318 4323 368 4357
rect 252 4316 304 4323
rect 316 4316 368 4323
rect 380 4316 432 4368
rect 444 4316 496 4368
rect 508 4357 560 4368
rect 508 4323 539 4357
rect 539 4323 560 4357
rect 508 4316 560 4323
rect 162 4309 171 4315
rect 171 4309 205 4315
rect 205 4309 214 4315
rect 162 4281 171 4292
rect 171 4281 205 4292
rect 205 4281 214 4292
rect 162 4241 214 4281
rect 252 4281 304 4294
rect 316 4281 368 4294
rect 252 4247 284 4281
rect 284 4247 304 4281
rect 316 4247 318 4281
rect 318 4247 368 4281
rect 252 4242 304 4247
rect 316 4242 368 4247
rect 380 4242 432 4294
rect 444 4242 496 4294
rect 508 4281 560 4294
rect 508 4247 539 4281
rect 539 4247 560 4281
rect 508 4242 560 4247
rect 162 4240 171 4241
rect 171 4240 205 4241
rect 205 4240 214 4241
rect 162 4207 171 4223
rect 171 4207 205 4223
rect 205 4207 214 4223
rect 162 4171 214 4207
rect 252 4205 304 4220
rect 316 4205 368 4220
rect 252 4171 284 4205
rect 284 4171 304 4205
rect 316 4171 318 4205
rect 318 4171 368 4205
rect 252 4168 304 4171
rect 316 4168 368 4171
rect 380 4168 432 4220
rect 444 4168 496 4220
rect 508 4205 560 4220
rect 508 4171 539 4205
rect 539 4171 560 4205
rect 508 4168 560 4171
rect 162 3245 171 3276
rect 171 3245 205 3276
rect 205 3245 214 3276
rect 162 3224 214 3245
rect 162 3205 214 3207
rect 162 3171 171 3205
rect 171 3171 205 3205
rect 205 3171 214 3205
rect 162 3155 214 3171
rect 162 3131 214 3138
rect 162 3097 171 3131
rect 171 3097 205 3131
rect 205 3097 214 3131
rect 162 3086 214 3097
rect 162 3057 214 3069
rect 162 3023 171 3057
rect 171 3023 205 3057
rect 205 3023 214 3057
rect 162 3017 214 3023
rect 167 2668 198 2702
rect 198 2668 219 2702
rect 167 2650 219 2668
rect 245 2668 266 2702
rect 266 2668 297 2702
rect 245 2650 297 2668
rect 167 2627 219 2635
rect 167 2593 198 2627
rect 198 2593 219 2627
rect 167 2583 219 2593
rect 245 2627 297 2635
rect 245 2593 266 2627
rect 266 2593 297 2627
rect 245 2583 297 2593
rect 167 2551 219 2568
rect 167 2517 198 2551
rect 198 2517 219 2551
rect 167 2516 219 2517
rect 245 2551 297 2568
rect 245 2517 266 2551
rect 266 2517 297 2551
rect 245 2516 297 2517
rect 167 2236 198 2270
rect 198 2236 219 2270
rect 167 2218 219 2236
rect 245 2236 266 2270
rect 266 2236 297 2270
rect 245 2218 297 2236
rect 167 2195 219 2203
rect 167 2161 198 2195
rect 198 2161 219 2195
rect 167 2151 219 2161
rect 245 2195 297 2203
rect 245 2161 266 2195
rect 266 2161 297 2195
rect 245 2151 297 2161
rect 167 2119 219 2136
rect 167 2085 198 2119
rect 198 2085 219 2119
rect 167 2084 219 2085
rect 245 2119 297 2136
rect 245 2085 266 2119
rect 266 2085 297 2119
rect 245 2084 297 2085
rect 160 1394 212 1409
rect 258 1399 310 1409
rect 160 1360 167 1394
rect 167 1360 201 1394
rect 201 1360 212 1394
rect 258 1365 289 1399
rect 289 1365 310 1399
rect 160 1357 212 1360
rect 258 1357 310 1365
rect 160 1320 212 1344
rect 258 1326 310 1344
rect 160 1292 167 1320
rect 167 1292 201 1320
rect 201 1292 212 1320
rect 258 1292 289 1326
rect 289 1292 310 1326
rect 160 1246 212 1279
rect 258 1253 310 1279
rect 160 1227 167 1246
rect 167 1227 201 1246
rect 201 1227 212 1246
rect 258 1227 289 1253
rect 289 1227 310 1253
rect 160 1212 167 1214
rect 167 1212 201 1214
rect 201 1212 212 1214
rect 160 1172 212 1212
rect 258 1180 310 1214
rect 160 1162 167 1172
rect 167 1162 201 1172
rect 201 1162 212 1172
rect 258 1162 289 1180
rect 289 1162 310 1180
rect 160 1138 167 1149
rect 167 1138 201 1149
rect 201 1138 212 1149
rect 258 1146 289 1149
rect 289 1146 310 1149
rect 160 1098 212 1138
rect 258 1107 310 1146
rect 160 1097 167 1098
rect 167 1097 201 1098
rect 201 1097 212 1098
rect 258 1097 289 1107
rect 289 1097 310 1107
rect 160 1064 167 1084
rect 167 1064 201 1084
rect 201 1064 212 1084
rect 258 1073 289 1084
rect 289 1073 310 1084
rect 160 1032 212 1064
rect 258 1034 310 1073
rect 258 1032 289 1034
rect 289 1032 310 1034
rect 160 991 167 1018
rect 167 991 201 1018
rect 201 991 212 1018
rect 258 1000 289 1018
rect 289 1000 310 1018
rect 160 966 212 991
rect 258 966 310 1000
rect 160 918 167 952
rect 167 918 201 952
rect 201 918 212 952
rect 258 927 289 952
rect 289 927 310 952
rect 160 900 212 918
rect 258 900 310 927
rect 160 879 212 886
rect 160 845 167 879
rect 167 845 201 879
rect 201 845 212 879
rect 258 854 289 886
rect 289 854 310 886
rect 160 834 212 845
rect 258 834 310 854
<< metal2 >>
rect 152 10292 310 10298
rect 152 10224 154 10292
rect 206 10280 258 10292
rect 310 10280 312 10289
rect 210 10224 256 10280
rect 152 10188 312 10224
rect 152 10121 154 10188
rect 206 10177 258 10188
rect 310 10177 312 10188
rect 210 10121 256 10177
rect 152 10083 312 10121
rect 152 10018 154 10083
rect 206 10074 258 10083
rect 310 10074 312 10083
rect 210 10018 256 10074
rect 152 9978 312 10018
rect 152 9915 154 9978
rect 206 9971 258 9978
rect 310 9971 312 9978
rect 210 9915 256 9971
rect 152 9873 312 9915
rect 152 9811 154 9873
rect 206 9867 258 9873
rect 310 9867 312 9873
rect 210 9811 256 9867
rect 152 9768 312 9811
rect 152 9707 154 9768
rect 206 9763 258 9768
rect 310 9763 312 9768
rect 210 9707 256 9763
rect 152 9698 312 9707
rect 152 8488 223 9698
rect 152 8479 312 8488
rect 152 8423 154 8479
rect 210 8423 256 8479
rect 152 8412 312 8423
rect 152 8295 154 8412
rect 206 8376 258 8412
rect 310 8376 312 8412
rect 210 8320 256 8376
rect 206 8295 258 8320
rect 310 8295 312 8320
rect 152 8282 312 8295
rect 152 8099 154 8282
rect 206 8273 258 8282
rect 310 8273 312 8282
rect 210 8217 256 8273
rect 206 8170 258 8217
rect 310 8170 312 8217
rect 210 8114 256 8170
rect 206 8099 258 8114
rect 310 8099 312 8114
rect 152 8085 312 8099
rect 152 7967 154 8085
rect 206 8066 258 8085
rect 310 8066 312 8085
rect 210 8010 256 8066
rect 206 7967 258 8010
rect 310 7967 312 8010
rect 152 7962 312 7967
rect 152 7901 154 7962
rect 210 7906 256 7962
rect 206 7901 258 7906
rect 310 7901 312 7906
rect 152 7897 312 7901
rect 152 7895 310 7897
rect 152 7087 223 7895
rect 152 7035 162 7087
rect 214 7035 223 7087
rect 152 7022 223 7035
rect 152 6970 162 7022
rect 214 6970 223 7022
rect 152 6957 223 6970
rect 152 6905 162 6957
rect 214 6905 223 6957
rect 152 6892 223 6905
rect 152 6840 162 6892
rect 214 6840 223 6892
rect 152 6833 223 6840
tri 223 6833 483 7093 sw
rect 152 6826 586 6833
rect 152 6774 162 6826
rect 214 6774 586 6826
rect 152 6760 586 6774
rect 152 6708 162 6760
rect 214 6708 586 6760
rect 152 6694 586 6708
rect 152 6672 162 6694
rect 214 6672 586 6694
rect 152 6616 154 6672
rect 214 6642 256 6672
rect 210 6628 256 6642
rect 214 6616 256 6628
rect 312 6616 586 6672
rect 152 6576 162 6616
rect 214 6576 586 6616
rect 152 6569 586 6576
rect 152 6513 154 6569
rect 210 6562 256 6569
rect 214 6513 256 6562
rect 312 6513 586 6569
rect 152 6510 162 6513
rect 214 6510 586 6513
rect 152 6496 586 6510
rect 152 6466 162 6496
rect 214 6466 586 6496
rect 152 6410 154 6466
rect 214 6444 256 6466
rect 210 6430 256 6444
rect 214 6410 256 6430
rect 312 6410 586 6466
rect 152 6378 162 6410
rect 214 6378 586 6410
rect 152 6364 586 6378
rect 152 6363 162 6364
rect 214 6363 586 6364
rect 152 6307 154 6363
rect 214 6312 256 6363
rect 210 6307 256 6312
rect 312 6307 586 6363
rect 152 6298 586 6307
rect 152 6259 162 6298
rect 214 6259 586 6298
rect 152 6203 154 6259
rect 214 6246 256 6259
rect 210 6232 256 6246
rect 214 6203 256 6232
rect 312 6203 586 6259
rect 152 6180 162 6203
rect 214 6180 586 6203
rect 152 6166 586 6180
rect 152 6155 162 6166
rect 214 6155 586 6166
rect 152 6099 154 6155
rect 214 6114 256 6155
rect 210 6100 256 6114
rect 214 6099 256 6100
rect 312 6099 586 6155
rect 152 6048 162 6099
rect 214 6071 586 6099
rect 214 6048 252 6071
rect 152 6034 252 6048
rect 152 5982 162 6034
rect 214 6019 252 6034
rect 304 6019 316 6071
rect 368 6019 380 6071
rect 432 6019 444 6071
rect 496 6019 508 6071
rect 560 6019 586 6071
rect 214 6002 586 6019
rect 214 5982 252 6002
rect 152 5968 252 5982
rect 152 5916 162 5968
rect 214 5950 252 5968
rect 304 5950 316 6002
rect 368 5950 380 6002
rect 432 5950 444 6002
rect 496 5950 508 6002
rect 560 5950 586 6002
rect 214 5933 586 5950
rect 214 5916 252 5933
rect 152 5902 252 5916
rect 152 5850 162 5902
rect 214 5881 252 5902
rect 304 5881 316 5933
rect 368 5881 380 5933
rect 432 5881 444 5933
rect 496 5881 508 5933
rect 560 5881 586 5933
rect 214 5864 586 5881
rect 214 5850 252 5864
rect 152 5836 252 5850
rect 152 5784 162 5836
rect 214 5812 252 5836
rect 304 5812 316 5864
rect 368 5812 380 5864
rect 432 5812 444 5864
rect 496 5812 508 5864
rect 560 5812 586 5864
rect 214 5795 586 5812
rect 214 5784 252 5795
rect 152 5770 252 5784
rect 152 5718 162 5770
rect 214 5743 252 5770
rect 304 5743 316 5795
rect 368 5743 380 5795
rect 432 5743 444 5795
rect 496 5743 508 5795
rect 560 5743 586 5795
rect 214 5726 586 5743
rect 214 5718 252 5726
rect 152 5704 252 5718
rect 152 5652 162 5704
rect 214 5674 252 5704
rect 304 5674 316 5726
rect 368 5674 380 5726
rect 432 5674 444 5726
rect 496 5674 508 5726
rect 560 5674 586 5726
rect 214 5657 586 5674
rect 214 5652 252 5657
rect 152 5638 252 5652
rect 152 5586 162 5638
rect 214 5605 252 5638
rect 304 5605 316 5657
rect 368 5605 380 5657
rect 432 5605 444 5657
rect 496 5605 508 5657
rect 560 5605 586 5657
rect 214 5588 586 5605
rect 214 5586 252 5588
rect 152 5572 252 5586
rect 152 5520 162 5572
rect 214 5536 252 5572
rect 304 5536 316 5588
rect 368 5536 380 5588
rect 432 5536 444 5588
rect 496 5536 508 5588
rect 560 5536 586 5588
rect 214 5520 586 5536
rect 152 5519 586 5520
rect 152 5506 252 5519
rect 152 5454 162 5506
rect 214 5467 252 5506
rect 304 5467 316 5519
rect 368 5467 380 5519
rect 432 5467 444 5519
rect 496 5467 508 5519
rect 560 5467 586 5519
rect 214 5454 586 5467
rect 152 5449 586 5454
rect 152 5440 252 5449
rect 152 5388 162 5440
rect 214 5397 252 5440
rect 304 5397 316 5449
rect 368 5397 380 5449
rect 432 5397 444 5449
rect 496 5397 508 5449
rect 560 5397 586 5449
rect 214 5388 586 5397
rect 152 5379 586 5388
rect 152 5374 252 5379
rect 152 5322 162 5374
rect 214 5327 252 5374
rect 304 5327 316 5379
rect 368 5327 380 5379
rect 432 5327 444 5379
rect 496 5327 508 5379
rect 560 5327 586 5379
rect 214 5322 586 5327
rect 152 5316 586 5322
rect 153 5031 319 5201
tri 319 5031 489 5201 sw
rect 153 4906 579 5031
rect 153 4868 162 4906
rect 214 4868 579 4906
rect 214 4854 263 4868
rect 209 4838 263 4854
rect 214 4812 263 4838
rect 319 4812 579 4868
rect 153 4786 162 4812
rect 214 4786 579 4812
rect 153 4770 579 4786
rect 153 4765 162 4770
rect 214 4765 579 4770
rect 214 4718 263 4765
rect 209 4709 263 4718
rect 319 4709 579 4765
rect 153 4702 579 4709
rect 153 4662 162 4702
rect 214 4664 579 4702
rect 214 4650 252 4664
rect 304 4662 316 4664
rect 209 4634 252 4650
rect 214 4612 252 4634
rect 368 4612 380 4664
rect 432 4612 444 4664
rect 496 4612 508 4664
rect 560 4612 579 4664
rect 214 4606 263 4612
rect 319 4606 579 4612
rect 153 4582 162 4606
rect 214 4590 579 4606
rect 214 4582 252 4590
rect 153 4566 252 4582
rect 153 4559 162 4566
rect 214 4538 252 4566
rect 304 4559 316 4590
rect 368 4538 380 4590
rect 432 4538 444 4590
rect 496 4538 508 4590
rect 560 4538 579 4590
rect 214 4516 263 4538
rect 319 4516 579 4538
rect 214 4514 252 4516
rect 209 4503 252 4514
rect 153 4498 252 4503
rect 153 4455 162 4498
rect 214 4464 252 4498
rect 304 4464 316 4503
rect 368 4464 380 4516
rect 432 4464 444 4516
rect 496 4464 508 4516
rect 560 4464 579 4516
rect 214 4455 579 4464
rect 214 4446 263 4455
rect 209 4442 263 4446
rect 319 4442 579 4455
rect 209 4430 252 4442
rect 153 4378 162 4399
rect 214 4390 252 4430
rect 304 4390 316 4399
rect 368 4390 380 4442
rect 432 4390 444 4442
rect 496 4390 508 4442
rect 560 4390 579 4442
rect 214 4378 579 4390
rect 153 4368 579 4378
rect 153 4361 252 4368
rect 153 4351 162 4361
rect 214 4316 252 4361
rect 304 4351 316 4368
rect 368 4316 380 4368
rect 432 4316 444 4368
rect 496 4316 508 4368
rect 560 4316 579 4368
rect 214 4309 263 4316
rect 209 4295 263 4309
rect 319 4295 579 4316
rect 153 4294 579 4295
rect 153 4292 252 4294
rect 153 4240 162 4292
rect 214 4242 252 4292
rect 304 4242 316 4294
rect 368 4242 380 4294
rect 432 4242 444 4294
rect 496 4242 508 4294
rect 560 4242 579 4294
rect 214 4240 579 4242
rect 153 4223 579 4240
rect 153 4171 162 4223
rect 214 4220 579 4223
rect 214 4171 252 4220
rect 153 4168 252 4171
rect 304 4168 316 4220
rect 368 4168 380 4220
rect 432 4168 444 4220
rect 496 4168 508 4220
rect 560 4168 579 4220
rect 153 4162 579 4168
rect 162 3276 311 3283
rect 214 3224 311 3276
rect 162 3207 311 3224
rect 214 3155 311 3207
rect 162 3138 311 3155
rect 214 3086 311 3138
rect 162 3069 311 3086
rect 214 3017 311 3069
rect 162 2702 311 3017
rect 162 2650 167 2702
rect 219 2650 245 2702
rect 297 2650 311 2702
rect 162 2635 311 2650
rect 162 2583 167 2635
rect 219 2583 245 2635
rect 297 2583 311 2635
rect 162 2568 311 2583
rect 162 2516 167 2568
rect 219 2516 245 2568
rect 297 2516 311 2568
rect 162 2270 311 2516
rect 162 2218 167 2270
rect 219 2218 245 2270
rect 297 2218 311 2270
rect 162 2203 311 2218
rect 162 2151 167 2203
rect 219 2151 245 2203
rect 297 2151 311 2203
rect 162 2136 311 2151
rect 162 2084 167 2136
rect 219 2084 245 2136
rect 297 2084 311 2136
rect 162 1579 311 2084
rect 162 1570 310 1579
rect 218 1514 254 1570
rect 162 1486 310 1514
rect 218 1430 254 1486
tri 160 1415 162 1417 se
rect 162 1415 310 1430
rect 160 1409 310 1415
rect 212 1402 258 1409
rect 160 1346 162 1357
rect 218 1346 254 1402
rect 160 1344 310 1346
rect 212 1318 258 1344
rect 160 1279 162 1292
rect 218 1262 254 1318
rect 212 1233 258 1262
rect 160 1214 162 1227
rect 218 1177 254 1233
rect 212 1162 258 1177
rect 160 1149 310 1162
rect 212 1148 258 1149
rect 160 1092 162 1097
rect 218 1092 254 1148
rect 160 1084 310 1092
rect 212 1063 258 1084
rect 160 1018 162 1032
rect 218 1007 254 1063
rect 212 966 258 1007
rect 160 952 310 966
rect 212 900 258 952
rect 160 886 310 900
rect 212 834 258 886
rect 160 828 310 834
<< via2 >>
rect 154 10240 206 10280
rect 206 10240 210 10280
rect 154 10224 210 10240
rect 256 10240 258 10280
rect 258 10240 310 10280
rect 310 10240 312 10280
rect 256 10224 312 10240
rect 154 10136 206 10177
rect 206 10136 210 10177
rect 154 10121 210 10136
rect 256 10136 258 10177
rect 258 10136 310 10177
rect 310 10136 312 10177
rect 256 10121 312 10136
rect 154 10031 206 10074
rect 206 10031 210 10074
rect 154 10018 210 10031
rect 256 10031 258 10074
rect 258 10031 310 10074
rect 310 10031 312 10074
rect 256 10018 312 10031
rect 154 9926 206 9971
rect 206 9926 210 9971
rect 154 9915 210 9926
rect 256 9926 258 9971
rect 258 9926 310 9971
rect 310 9926 312 9971
rect 256 9915 312 9926
rect 154 9821 206 9867
rect 206 9821 210 9867
rect 154 9811 210 9821
rect 256 9821 258 9867
rect 258 9821 310 9867
rect 310 9821 312 9867
rect 256 9811 312 9821
rect 154 9716 206 9763
rect 206 9716 210 9763
rect 154 9707 210 9716
rect 256 9716 258 9763
rect 258 9716 310 9763
rect 310 9716 312 9763
rect 256 9707 312 9716
rect 154 8477 210 8479
rect 154 8425 206 8477
rect 206 8425 210 8477
rect 154 8423 210 8425
rect 256 8477 312 8479
rect 256 8425 258 8477
rect 258 8425 310 8477
rect 310 8425 312 8477
rect 256 8423 312 8425
rect 154 8360 206 8376
rect 206 8360 210 8376
rect 154 8347 210 8360
rect 154 8320 206 8347
rect 206 8320 210 8347
rect 256 8360 258 8376
rect 258 8360 310 8376
rect 310 8360 312 8376
rect 256 8347 312 8360
rect 256 8320 258 8347
rect 258 8320 310 8347
rect 310 8320 312 8347
rect 154 8230 206 8273
rect 206 8230 210 8273
rect 154 8217 210 8230
rect 256 8230 258 8273
rect 258 8230 310 8273
rect 310 8230 312 8273
rect 256 8217 312 8230
rect 154 8165 206 8170
rect 206 8165 210 8170
rect 154 8151 210 8165
rect 154 8114 206 8151
rect 206 8114 210 8151
rect 256 8165 258 8170
rect 258 8165 310 8170
rect 310 8165 312 8170
rect 256 8151 312 8165
rect 256 8114 258 8151
rect 258 8114 310 8151
rect 310 8114 312 8151
rect 154 8033 206 8066
rect 206 8033 210 8066
rect 154 8019 210 8033
rect 154 8010 206 8019
rect 206 8010 210 8019
rect 256 8033 258 8066
rect 258 8033 310 8066
rect 310 8033 312 8066
rect 256 8019 312 8033
rect 256 8010 258 8019
rect 258 8010 310 8019
rect 310 8010 312 8019
rect 154 7953 210 7962
rect 154 7906 206 7953
rect 206 7906 210 7953
rect 256 7953 312 7962
rect 256 7906 258 7953
rect 258 7906 310 7953
rect 310 7906 312 7953
rect 154 6642 162 6672
rect 162 6642 210 6672
rect 154 6628 210 6642
rect 154 6616 162 6628
rect 162 6616 210 6628
rect 256 6616 312 6672
rect 154 6562 210 6569
rect 154 6513 162 6562
rect 162 6513 210 6562
rect 256 6513 312 6569
rect 154 6444 162 6466
rect 162 6444 210 6466
rect 154 6430 210 6444
rect 154 6410 162 6430
rect 162 6410 210 6430
rect 256 6410 312 6466
rect 154 6312 162 6363
rect 162 6312 210 6363
rect 154 6307 210 6312
rect 256 6307 312 6363
rect 154 6246 162 6259
rect 162 6246 210 6259
rect 154 6232 210 6246
rect 154 6203 162 6232
rect 162 6203 210 6232
rect 256 6203 312 6259
rect 154 6114 162 6155
rect 162 6114 210 6155
rect 154 6100 210 6114
rect 154 6099 162 6100
rect 162 6099 210 6100
rect 256 6099 312 6155
rect 153 4854 162 4868
rect 162 4854 209 4868
rect 153 4838 209 4854
rect 153 4812 162 4838
rect 162 4812 209 4838
rect 263 4812 319 4868
rect 153 4718 162 4765
rect 162 4718 209 4765
rect 153 4709 209 4718
rect 263 4709 319 4765
rect 153 4650 162 4662
rect 162 4650 209 4662
rect 153 4634 209 4650
rect 153 4606 162 4634
rect 162 4606 209 4634
rect 263 4612 304 4662
rect 304 4612 316 4662
rect 316 4612 319 4662
rect 263 4606 319 4612
rect 153 4514 162 4559
rect 162 4514 209 4559
rect 263 4538 304 4559
rect 304 4538 316 4559
rect 316 4538 319 4559
rect 263 4516 319 4538
rect 153 4503 209 4514
rect 263 4503 304 4516
rect 304 4503 316 4516
rect 316 4503 319 4516
rect 153 4446 162 4455
rect 162 4446 209 4455
rect 153 4430 209 4446
rect 263 4442 319 4455
rect 153 4399 162 4430
rect 162 4399 209 4430
rect 263 4399 304 4442
rect 304 4399 316 4442
rect 316 4399 319 4442
rect 153 4309 162 4351
rect 162 4309 209 4351
rect 263 4316 304 4351
rect 304 4316 316 4351
rect 316 4316 319 4351
rect 153 4295 209 4309
rect 263 4295 319 4316
rect 162 1514 218 1570
rect 254 1514 310 1570
rect 162 1430 218 1486
rect 254 1430 310 1486
rect 162 1357 212 1402
rect 212 1357 218 1402
rect 162 1346 218 1357
rect 254 1357 258 1402
rect 258 1357 310 1402
rect 254 1346 310 1357
rect 162 1292 212 1318
rect 212 1292 218 1318
rect 162 1279 218 1292
rect 162 1262 212 1279
rect 212 1262 218 1279
rect 254 1292 258 1318
rect 258 1292 310 1318
rect 254 1279 310 1292
rect 254 1262 258 1279
rect 258 1262 310 1279
rect 162 1227 212 1233
rect 212 1227 218 1233
rect 162 1214 218 1227
rect 162 1177 212 1214
rect 212 1177 218 1214
rect 254 1227 258 1233
rect 258 1227 310 1233
rect 254 1214 310 1227
rect 254 1177 258 1214
rect 258 1177 310 1214
rect 162 1097 212 1148
rect 212 1097 218 1148
rect 162 1092 218 1097
rect 254 1097 258 1148
rect 258 1097 310 1148
rect 254 1092 310 1097
rect 162 1032 212 1063
rect 212 1032 218 1063
rect 162 1018 218 1032
rect 162 1007 212 1018
rect 212 1007 218 1018
rect 254 1032 258 1063
rect 258 1032 310 1063
rect 254 1018 310 1032
rect 254 1007 258 1018
rect 258 1007 310 1018
<< metal3 >>
rect 149 10280 317 10285
rect 149 10224 154 10280
rect 210 10224 256 10280
rect 312 10224 317 10280
rect 149 10177 317 10224
rect 149 10121 154 10177
rect 210 10121 256 10177
rect 312 10121 317 10177
rect 149 10074 317 10121
rect 149 10018 154 10074
rect 210 10018 256 10074
rect 312 10018 317 10074
rect 149 9971 317 10018
rect 149 9915 154 9971
rect 210 9915 256 9971
rect 312 9915 317 9971
rect 149 9867 317 9915
rect 149 9811 154 9867
rect 210 9811 256 9867
rect 312 9811 317 9867
rect 149 9763 317 9811
rect 149 9707 154 9763
rect 210 9707 256 9763
rect 312 9707 317 9763
rect 149 9702 317 9707
rect 149 8479 317 8484
rect 149 8423 154 8479
rect 210 8423 256 8479
rect 312 8423 317 8479
rect 149 8376 317 8423
rect 149 8320 154 8376
rect 210 8320 256 8376
rect 312 8320 317 8376
rect 149 8273 317 8320
rect 149 8217 154 8273
rect 210 8217 256 8273
rect 312 8217 317 8273
rect 149 8170 317 8217
rect 149 8114 154 8170
rect 210 8114 256 8170
rect 312 8114 317 8170
rect 149 8066 317 8114
rect 149 8010 154 8066
rect 210 8010 256 8066
rect 312 8010 317 8066
rect 149 7962 317 8010
rect 149 7906 154 7962
rect 210 7906 256 7962
rect 312 7906 317 7962
rect 149 7901 317 7906
rect 149 6672 317 6677
rect 149 6616 154 6672
rect 210 6616 256 6672
rect 312 6616 317 6672
rect 149 6569 317 6616
rect 149 6513 154 6569
rect 210 6513 256 6569
rect 312 6513 317 6569
rect 149 6466 317 6513
rect 149 6410 154 6466
rect 210 6410 256 6466
rect 312 6410 317 6466
rect 149 6363 317 6410
rect 149 6307 154 6363
rect 210 6307 256 6363
rect 312 6307 317 6363
rect 149 6259 317 6307
rect 149 6203 154 6259
rect 210 6203 256 6259
rect 312 6203 317 6259
rect 149 6155 317 6203
rect 149 6099 154 6155
rect 210 6099 256 6155
rect 312 6099 317 6155
rect 149 6094 317 6099
rect 148 4868 324 4873
rect 148 4812 153 4868
rect 209 4812 263 4868
rect 319 4812 324 4868
rect 148 4765 324 4812
rect 148 4709 153 4765
rect 209 4709 263 4765
rect 319 4709 324 4765
rect 148 4662 324 4709
rect 148 4606 153 4662
rect 209 4606 263 4662
rect 319 4606 324 4662
rect 148 4559 324 4606
rect 148 4503 153 4559
rect 209 4503 263 4559
rect 319 4503 324 4559
rect 148 4455 324 4503
rect 148 4399 153 4455
rect 209 4399 263 4455
rect 319 4399 324 4455
rect 148 4351 324 4399
rect 148 4295 153 4351
rect 209 4295 263 4351
rect 319 4295 324 4351
rect 148 4290 324 4295
rect 157 1570 315 1575
rect 157 1514 162 1570
rect 218 1514 254 1570
rect 310 1514 315 1570
rect 157 1486 315 1514
rect 157 1430 162 1486
rect 218 1430 254 1486
rect 310 1430 315 1486
rect 157 1402 315 1430
rect 157 1346 162 1402
rect 218 1346 254 1402
rect 310 1346 315 1402
rect 157 1318 315 1346
rect 157 1262 162 1318
rect 218 1262 254 1318
rect 310 1262 315 1318
rect 157 1233 315 1262
rect 157 1177 162 1233
rect 218 1177 254 1233
rect 310 1177 315 1233
rect 157 1148 315 1177
rect 157 1092 162 1148
rect 218 1092 254 1148
rect 310 1092 315 1148
rect 157 1063 315 1092
rect 157 1007 162 1063
rect 218 1007 254 1063
rect 310 1007 315 1063
rect 157 1002 315 1007
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_0
timestamp 1679235063
transform 1 0 415 0 -1 3593
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_1
timestamp 1679235063
transform 1 0 415 0 -1 4714
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_2
timestamp 1679235063
transform 1 0 415 0 -1 2472
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_5595914180850  sky130_fd_pr__nfet_01v8__example_5595914180850_3
timestamp 1679235063
transform 1 0 415 0 1 362
box -1 0 121 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_0
timestamp 1679235063
transform 1 0 456 0 1 1384
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_1
timestamp 1679235063
transform 1 0 456 0 1 2503
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180839  sky130_fd_pr__via_pol1__example_5595914180839_2
timestamp 1679235063
transform 1 0 456 0 1 3624
box 0 0 1 1
<< labels >>
flabel comment s 212 3515 212 3515 0 FreeSans 400 90 0 0 CONDIODE
flabel metal1 s 124 2328 176 2458 0 FreeSans 200 0 0 0 PD_H
port 2 nsew
flabel metal1 s -50 1898 0 2028 0 FreeSans 200 0 0 0 PAD
port 3 nsew
flabel metal1 s -50 2758 0 2888 0 FreeSans 200 0 0 0 PAD
port 3 nsew
<< properties >>
string GDS_END 43449484
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43338452
<< end >>
