magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 1 21 1597 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 419 47 449 177
rect 503 47 533 177
rect 791 47 821 177
rect 875 47 905 177
rect 959 47 989 177
rect 1049 47 1079 177
rect 1237 47 1267 177
rect 1321 47 1351 177
rect 1405 47 1435 177
rect 1489 47 1519 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 519 297 549 497
rect 603 297 633 497
rect 791 297 821 497
rect 875 297 905 497
rect 959 297 989 497
rect 1049 297 1079 497
rect 1237 297 1267 497
rect 1321 297 1351 497
rect 1405 297 1435 497
rect 1489 297 1519 497
<< ndiff >>
rect 27 118 79 177
rect 27 84 35 118
rect 69 84 79 118
rect 27 47 79 84
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 161 247 177
rect 193 127 203 161
rect 237 127 247 161
rect 193 47 247 127
rect 277 93 331 177
rect 277 59 287 93
rect 321 59 331 93
rect 277 47 331 59
rect 361 161 419 177
rect 361 127 375 161
rect 409 127 419 161
rect 361 47 419 127
rect 449 93 503 177
rect 449 59 459 93
rect 493 59 503 93
rect 449 47 503 59
rect 533 118 585 177
rect 533 84 543 118
rect 577 84 585 118
rect 533 47 585 84
rect 739 161 791 177
rect 739 127 747 161
rect 781 127 791 161
rect 739 47 791 127
rect 821 93 875 177
rect 821 59 831 93
rect 865 59 875 93
rect 821 47 875 59
rect 905 161 959 177
rect 905 127 915 161
rect 949 127 959 161
rect 905 47 959 127
rect 989 93 1049 177
rect 989 59 1005 93
rect 1039 59 1049 93
rect 989 47 1049 59
rect 1079 161 1131 177
rect 1079 127 1089 161
rect 1123 127 1131 161
rect 1079 47 1131 127
rect 1185 161 1237 177
rect 1185 127 1193 161
rect 1227 127 1237 161
rect 1185 93 1237 127
rect 1185 59 1193 93
rect 1227 59 1237 93
rect 1185 47 1237 59
rect 1267 161 1321 177
rect 1267 127 1277 161
rect 1311 127 1321 161
rect 1267 93 1321 127
rect 1267 59 1277 93
rect 1311 59 1321 93
rect 1267 47 1321 59
rect 1351 93 1405 177
rect 1351 59 1361 93
rect 1395 59 1405 93
rect 1351 47 1405 59
rect 1435 161 1489 177
rect 1435 127 1445 161
rect 1479 127 1489 161
rect 1435 93 1489 127
rect 1435 59 1445 93
rect 1479 59 1489 93
rect 1435 47 1489 59
rect 1519 93 1571 177
rect 1519 59 1529 93
rect 1563 59 1571 93
rect 1519 47 1571 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 297 163 383
rect 193 485 247 497
rect 193 451 203 485
rect 237 451 247 485
rect 193 417 247 451
rect 193 383 203 417
rect 237 383 247 417
rect 193 349 247 383
rect 193 315 203 349
rect 237 315 247 349
rect 193 297 247 315
rect 277 390 331 497
rect 277 356 287 390
rect 321 356 331 390
rect 277 297 331 356
rect 361 485 413 497
rect 361 451 371 485
rect 405 451 413 485
rect 361 417 413 451
rect 361 383 371 417
rect 405 383 413 417
rect 361 297 413 383
rect 467 485 519 497
rect 467 451 475 485
rect 509 451 519 485
rect 467 417 519 451
rect 467 383 475 417
rect 509 383 519 417
rect 467 349 519 383
rect 467 315 475 349
rect 509 315 519 349
rect 467 297 519 315
rect 549 390 603 497
rect 549 356 559 390
rect 593 356 603 390
rect 549 297 603 356
rect 633 485 685 497
rect 633 451 643 485
rect 677 451 685 485
rect 633 417 685 451
rect 633 383 643 417
rect 677 383 685 417
rect 633 349 685 383
rect 633 315 643 349
rect 677 315 685 349
rect 633 297 685 315
rect 739 485 791 497
rect 739 451 747 485
rect 781 451 791 485
rect 739 417 791 451
rect 739 383 747 417
rect 781 383 791 417
rect 739 349 791 383
rect 739 315 747 349
rect 781 315 791 349
rect 739 297 791 315
rect 821 475 875 497
rect 821 441 831 475
rect 865 441 875 475
rect 821 297 875 441
rect 905 485 959 497
rect 905 451 915 485
rect 949 451 959 485
rect 905 417 959 451
rect 905 383 915 417
rect 949 383 959 417
rect 905 297 959 383
rect 989 407 1049 497
rect 989 373 1005 407
rect 1039 373 1049 407
rect 989 297 1049 373
rect 1079 485 1131 497
rect 1079 451 1089 485
rect 1123 451 1131 485
rect 1079 417 1131 451
rect 1079 383 1089 417
rect 1123 383 1131 417
rect 1079 349 1131 383
rect 1079 315 1089 349
rect 1123 315 1131 349
rect 1079 297 1131 315
rect 1185 485 1237 497
rect 1185 451 1193 485
rect 1227 451 1237 485
rect 1185 417 1237 451
rect 1185 383 1193 417
rect 1227 383 1237 417
rect 1185 297 1237 383
rect 1267 485 1321 497
rect 1267 451 1277 485
rect 1311 451 1321 485
rect 1267 417 1321 451
rect 1267 383 1277 417
rect 1311 383 1321 417
rect 1267 349 1321 383
rect 1267 315 1277 349
rect 1311 315 1321 349
rect 1267 297 1321 315
rect 1351 485 1405 497
rect 1351 451 1361 485
rect 1395 451 1405 485
rect 1351 417 1405 451
rect 1351 383 1361 417
rect 1395 383 1405 417
rect 1351 297 1405 383
rect 1435 485 1489 497
rect 1435 451 1445 485
rect 1479 451 1489 485
rect 1435 417 1489 451
rect 1435 383 1445 417
rect 1479 383 1489 417
rect 1435 349 1489 383
rect 1435 315 1445 349
rect 1479 315 1489 349
rect 1435 297 1489 315
rect 1519 485 1571 497
rect 1519 451 1529 485
rect 1563 451 1571 485
rect 1519 417 1571 451
rect 1519 383 1529 417
rect 1563 383 1571 417
rect 1519 297 1571 383
<< ndiffc >>
rect 35 84 69 118
rect 119 59 153 93
rect 203 127 237 161
rect 287 59 321 93
rect 375 127 409 161
rect 459 59 493 93
rect 543 84 577 118
rect 747 127 781 161
rect 831 59 865 93
rect 915 127 949 161
rect 1005 59 1039 93
rect 1089 127 1123 161
rect 1193 127 1227 161
rect 1193 59 1227 93
rect 1277 127 1311 161
rect 1277 59 1311 93
rect 1361 59 1395 93
rect 1445 127 1479 161
rect 1445 59 1479 93
rect 1529 59 1563 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 203 451 237 485
rect 203 383 237 417
rect 203 315 237 349
rect 287 356 321 390
rect 371 451 405 485
rect 371 383 405 417
rect 475 451 509 485
rect 475 383 509 417
rect 475 315 509 349
rect 559 356 593 390
rect 643 451 677 485
rect 643 383 677 417
rect 643 315 677 349
rect 747 451 781 485
rect 747 383 781 417
rect 747 315 781 349
rect 831 441 865 475
rect 915 451 949 485
rect 915 383 949 417
rect 1005 373 1039 407
rect 1089 451 1123 485
rect 1089 383 1123 417
rect 1089 315 1123 349
rect 1193 451 1227 485
rect 1193 383 1227 417
rect 1277 451 1311 485
rect 1277 383 1311 417
rect 1277 315 1311 349
rect 1361 451 1395 485
rect 1361 383 1395 417
rect 1445 451 1479 485
rect 1445 383 1479 417
rect 1445 315 1479 349
rect 1529 451 1563 485
rect 1529 383 1563 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 519 497 549 523
rect 603 497 633 523
rect 791 497 821 523
rect 875 497 905 523
rect 959 497 989 523
rect 1049 497 1079 523
rect 1237 497 1267 523
rect 1321 497 1351 523
rect 1405 497 1435 523
rect 1489 497 1519 523
rect 79 259 109 297
rect 163 259 193 297
rect 21 249 193 259
rect 21 215 76 249
rect 110 215 193 249
rect 21 205 193 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 259 277 297
rect 331 259 361 297
rect 519 259 549 297
rect 603 259 633 297
rect 791 259 821 297
rect 875 259 905 297
rect 247 249 361 259
rect 247 215 290 249
rect 324 215 361 249
rect 247 205 361 215
rect 247 177 277 205
rect 331 177 361 205
rect 419 249 633 259
rect 419 215 435 249
rect 469 215 633 249
rect 419 205 633 215
rect 780 249 905 259
rect 780 215 796 249
rect 830 215 905 249
rect 780 205 905 215
rect 419 177 449 205
rect 503 177 533 205
rect 791 177 821 205
rect 875 177 905 205
rect 959 259 989 297
rect 1049 259 1079 297
rect 1237 259 1267 297
rect 1321 259 1351 297
rect 1405 259 1435 297
rect 1489 259 1519 297
rect 959 249 1079 259
rect 959 215 1002 249
rect 1036 215 1079 249
rect 959 205 1079 215
rect 1178 249 1519 259
rect 1178 215 1194 249
rect 1228 215 1277 249
rect 1311 215 1361 249
rect 1395 215 1445 249
rect 1479 215 1519 249
rect 1178 205 1519 215
rect 959 177 989 205
rect 1049 177 1079 205
rect 1237 177 1267 205
rect 1321 177 1351 205
rect 1405 177 1435 205
rect 1489 177 1519 205
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 419 21 449 47
rect 503 21 533 47
rect 791 21 821 47
rect 875 21 905 47
rect 959 21 989 47
rect 1049 21 1079 47
rect 1237 21 1267 47
rect 1321 21 1351 47
rect 1405 21 1435 47
rect 1489 21 1519 47
<< polycont >>
rect 76 215 110 249
rect 290 215 324 249
rect 435 215 469 249
rect 796 215 830 249
rect 1002 215 1036 249
rect 1194 215 1228 249
rect 1277 215 1311 249
rect 1361 215 1395 249
rect 1445 215 1479 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 485 85 493
rect 17 451 35 485
rect 69 451 85 485
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 119 485 153 527
rect 119 417 153 451
rect 119 367 153 383
rect 187 485 421 493
rect 187 451 203 485
rect 237 459 371 485
rect 237 451 253 459
rect 187 417 253 451
rect 187 383 203 417
rect 237 383 253 417
rect 355 451 371 459
rect 405 451 421 485
rect 355 417 421 451
rect 17 315 35 349
rect 69 333 85 349
rect 187 349 253 383
rect 187 333 203 349
rect 69 315 203 333
rect 237 315 253 349
rect 17 289 253 315
rect 287 390 321 409
rect 355 383 371 417
rect 405 383 421 417
rect 355 372 421 383
rect 459 485 693 493
rect 459 451 475 485
rect 509 459 643 485
rect 509 451 525 459
rect 459 417 525 451
rect 459 383 475 417
rect 509 383 525 417
rect 627 451 643 459
rect 677 451 693 485
rect 627 417 693 451
rect 287 338 321 356
rect 459 349 525 383
rect 459 338 475 349
rect 287 315 475 338
rect 509 315 525 349
rect 287 289 525 315
rect 559 390 593 409
rect 559 255 593 356
rect 627 383 643 417
rect 677 383 693 417
rect 627 349 693 383
rect 627 315 643 349
rect 677 315 693 349
rect 627 289 693 315
rect 731 485 797 493
rect 731 451 747 485
rect 781 451 797 485
rect 731 417 797 451
rect 831 475 865 527
rect 831 425 865 441
rect 899 485 1139 493
rect 899 451 915 485
rect 949 457 1089 485
rect 949 451 965 457
rect 731 383 747 417
rect 781 391 797 417
rect 899 417 965 451
rect 1073 451 1089 457
rect 1123 451 1139 485
rect 899 391 915 417
rect 781 383 915 391
rect 949 383 965 417
rect 731 357 965 383
rect 1005 407 1039 423
rect 731 349 797 357
rect 731 315 747 349
rect 781 315 797 349
rect 1005 323 1039 373
rect 731 289 797 315
rect 880 289 1039 323
rect 1073 417 1139 451
rect 1073 383 1089 417
rect 1123 383 1139 417
rect 1073 349 1139 383
rect 1193 485 1227 527
rect 1193 417 1227 451
rect 1193 367 1227 383
rect 1261 485 1327 493
rect 1261 451 1277 485
rect 1311 451 1327 485
rect 1261 417 1327 451
rect 1261 383 1277 417
rect 1311 383 1327 417
rect 1073 315 1089 349
rect 1123 315 1139 349
rect 1073 289 1139 315
rect 1261 349 1327 383
rect 1361 485 1395 527
rect 1361 417 1395 451
rect 1361 367 1395 383
rect 1429 485 1495 493
rect 1429 451 1445 485
rect 1479 451 1495 485
rect 1429 417 1495 451
rect 1429 383 1445 417
rect 1479 383 1495 417
rect 1261 315 1277 349
rect 1311 333 1327 349
rect 1429 349 1495 383
rect 1529 485 1580 527
rect 1563 451 1580 485
rect 1529 417 1580 451
rect 1563 383 1580 417
rect 1529 367 1580 383
rect 1429 333 1445 349
rect 1311 315 1445 333
rect 1479 333 1495 349
rect 1479 315 1627 333
rect 1261 299 1627 315
rect 30 249 156 255
rect 30 215 76 249
rect 110 215 156 249
rect 214 249 340 255
rect 214 215 290 249
rect 324 215 340 249
rect 402 249 525 255
rect 402 215 435 249
rect 469 215 525 249
rect 559 221 729 255
rect 17 161 593 177
rect 17 127 203 161
rect 237 127 375 161
rect 409 127 593 161
rect 691 161 729 221
rect 774 249 846 255
rect 774 215 796 249
rect 830 215 846 249
rect 880 161 924 289
rect 958 249 1052 255
rect 958 215 1002 249
rect 1036 215 1052 249
rect 1104 249 1227 253
rect 1104 215 1194 249
rect 1228 215 1277 249
rect 1311 215 1361 249
rect 1395 215 1445 249
rect 1479 215 1495 249
rect 1104 161 1155 215
rect 1529 181 1627 299
rect 691 127 747 161
rect 781 127 915 161
rect 949 127 1089 161
rect 1123 127 1155 161
rect 1193 161 1227 177
rect 17 118 69 127
rect 17 84 35 118
rect 543 118 593 127
rect 17 51 69 84
rect 103 59 119 93
rect 153 59 287 93
rect 321 59 459 93
rect 493 59 509 93
rect 103 17 509 59
rect 577 93 593 118
rect 1193 93 1227 127
rect 577 84 831 93
rect 543 59 831 84
rect 865 59 1005 93
rect 1039 59 1139 93
rect 543 51 1139 59
rect 1193 17 1227 59
rect 1261 161 1627 181
rect 1261 127 1277 161
rect 1311 143 1445 161
rect 1311 127 1327 143
rect 1261 93 1327 127
rect 1429 127 1445 143
rect 1479 143 1627 161
rect 1479 127 1495 143
rect 1261 59 1277 93
rect 1311 59 1327 93
rect 1261 51 1327 59
rect 1361 93 1395 109
rect 1361 17 1395 59
rect 1429 93 1495 127
rect 1429 59 1445 93
rect 1479 59 1495 93
rect 1429 51 1495 59
rect 1529 93 1580 109
rect 1563 59 1580 93
rect 1529 17 1580 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 1593 153 1627 187 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 1593 221 1627 255 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 1593 289 1627 323 0 FreeSans 200 0 0 0 X
port 10 nsew signal output
flabel locali s 958 221 992 255 0 FreeSans 200 0 0 0 B2
port 5 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 774 221 808 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o32a_4
rlabel metal1 s 0 -48 1656 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 1480874
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1468626
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 8.280 0.000 
<< end >>
