magic
tech sky130A
magscale 1 2
timestamp 1679235063
use sky130_fd_io__tk_em1o_cdns_5595914180879  sky130_fd_io__tk_em1o_cdns_5595914180879_0
timestamp 1679235063
transform -1 0 15232 0 1 3026
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_55959141808327  sky130_fd_io__tk_em1o_cdns_55959141808327_0
timestamp 1679235063
transform -1 0 13342 0 1 3470
box 0 0 1 1
use sky130_fd_io__tk_em1o_cdns_55959141808328  sky130_fd_io__tk_em1o_cdns_55959141808328_0
timestamp 1679235063
transform 0 -1 12023 -1 0 4792
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180881  sky130_fd_io__tk_em1s_cdns_5595914180881_0
timestamp 1679235063
transform 1 0 16744 0 1 3552
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_0
timestamp 1679235063
transform 1 0 11787 0 1 4381
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180882  sky130_fd_io__tk_em1s_cdns_5595914180882_1
timestamp 1679235063
transform 1 0 11628 0 1 3386
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_0
timestamp 1679235063
transform 0 -1 12686 1 0 4032
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_55959141808288  sky130_fd_io__tk_em1s_cdns_55959141808288_1
timestamp 1679235063
transform 0 -1 13002 1 0 3881
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808134  sky130_fd_pr__nfet_01v8__example_55959141808134_0
timestamp 1679235063
transform -1 0 12901 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808304  sky130_fd_pr__nfet_01v8__example_55959141808304_0
timestamp 1679235063
transform 0 -1 12060 -1 0 4784
box -1 0 101 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_0
timestamp 1679235063
transform 1 0 13309 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_1
timestamp 1679235063
transform -1 0 13253 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_2
timestamp 1679235063
transform 1 0 12957 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808329  sky130_fd_pr__nfet_01v8__example_55959141808329_3
timestamp 1679235063
transform 1 0 12605 0 1 4311
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808330  sky130_fd_pr__nfet_01v8__example_55959141808330_0
timestamp 1679235063
transform -1 0 12293 0 1 4573
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808330  sky130_fd_pr__nfet_01v8__example_55959141808330_1
timestamp 1679235063
transform 0 1 12406 -1 0 4804
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808331  sky130_fd_pr__nfet_01v8__example_55959141808331_0
timestamp 1679235063
transform 1 0 11581 0 1 4311
box -1 0 457 1
use sky130_fd_pr__nfet_01v8__example_55959141808332  sky130_fd_pr__nfet_01v8__example_55959141808332_0
timestamp 1679235063
transform 1 0 12093 0 1 4311
box -1 0 457 1
use sky130_fd_pr__nfet_01v8__example_55959141808333  sky130_fd_pr__nfet_01v8__example_55959141808333_0
timestamp 1679235063
transform 0 -1 12662 1 0 3225
box -1 0 801 1
use sky130_fd_pr__nfet_01v8__example_55959141808334  sky130_fd_pr__nfet_01v8__example_55959141808334_0
timestamp 1679235063
transform 0 -1 12518 -1 0 4025
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808343  sky130_fd_pr__pfet_01v8__example_55959141808343_0
timestamp 1679235063
transform -1 0 17991 0 -1 4078
box -1 0 1193 1
use sky130_fd_pr__pfet_01v8__example_55959141808343  sky130_fd_pr__pfet_01v8__example_55959141808343_1
timestamp 1679235063
transform 1 0 13911 0 -1 4078
box -1 0 1193 1
use sky130_fd_pr__pfet_01v8__example_55959141808343  sky130_fd_pr__pfet_01v8__example_55959141808343_2
timestamp 1679235063
transform 1 0 15355 0 -1 4028
box -1 0 1193 1
use sky130_fd_pr__pfet_01v8__example_55959141808344  sky130_fd_pr__pfet_01v8__example_55959141808344_0
timestamp 1679235063
transform -1 0 19701 0 -1 4078
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808344  sky130_fd_pr__pfet_01v8__example_55959141808344_1
timestamp 1679235063
transform 1 0 19757 0 -1 4078
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808344  sky130_fd_pr__pfet_01v8__example_55959141808344_2
timestamp 1679235063
transform -1 0 13855 0 -1 4078
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808345  sky130_fd_pr__pfet_01v8__example_55959141808345_0
timestamp 1679235063
transform 0 -1 12990 1 0 3225
box -1 0 801 1
use sky130_fd_pr__pfet_01v8__example_55959141808346  sky130_fd_pr__pfet_01v8__example_55959141808346_0
timestamp 1679235063
transform 1 0 18867 0 -1 4078
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808346  sky130_fd_pr__pfet_01v8__example_55959141808346_1
timestamp 1679235063
transform 1 0 18243 0 -1 4078
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808347  sky130_fd_pr__pfet_01v8__example_55959141808347_0
timestamp 1679235063
transform -1 0 13503 0 -1 4073
box -1 0 257 1
use sky130_fd_pr__pfet_01v8__example_55959141808348  sky130_fd_pr__pfet_01v8__example_55959141808348_0
timestamp 1679235063
transform 1 0 17679 0 -1 4256
box -1 0 1601 1
use sky130_fd_pr__pfet_01v8__example_55959141808639  sky130_fd_pr__pfet_01v8__example_55959141808639_0
timestamp 1679235063
transform 1 0 13119 0 -1 3678
box -1 0 0 1
use sky130_fd_pr__pfet_01v8__example_55959141808640  sky130_fd_pr__pfet_01v8__example_55959141808640_0
timestamp 1679235063
transform 1 0 13261 0 -1 3678
box 0 0 1 1
use sky130_fd_pr__pfet_01v8__example_55959141808641  sky130_fd_pr__pfet_01v8__example_55959141808641_0
timestamp 1679235063
transform 1 0 13403 0 -1 3678
box 100 0 101 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1679235063
transform -1 0 13392 0 -1 3976
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1679235063
transform 1 0 12299 0 -1 3429
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1679235063
transform -1 0 12674 0 1 4036
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1679235063
transform 1 0 12990 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1679235063
transform -1 0 12736 0 1 4571
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1679235063
transform -1 0 13510 0 1 3030
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1679235063
transform 1 0 11718 0 1 4391
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1679235063
transform 1 0 12232 0 1 4387
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1679235063
transform 1 0 16368 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_9
timestamp 1679235063
transform 1 0 16056 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_10
timestamp 1679235063
transform 1 0 15744 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_11
timestamp 1679235063
transform 1 0 15432 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_12
timestamp 1679235063
transform 1 0 19796 0 1 3862
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_13
timestamp 1679235063
transform 0 1 13710 1 0 3868
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_14
timestamp 1679235063
transform -1 0 12990 0 -1 4013
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_15
timestamp 1679235063
transform 1 0 12056 0 1 4553
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_16
timestamp 1679235063
transform 1 0 13084 0 -1 3064
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_17
timestamp 1679235063
transform 1 0 13475 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_18
timestamp 1679235063
transform 1 0 13148 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_19
timestamp 1679235063
transform 1 0 17494 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_20
timestamp 1679235063
transform 1 0 17812 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_21
timestamp 1679235063
transform 1 0 16877 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_22
timestamp 1679235063
transform 1 0 17188 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_23
timestamp 1679235063
transform 1 0 15901 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_24
timestamp 1679235063
transform 1 0 16213 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_25
timestamp 1679235063
transform 1 0 16487 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_26
timestamp 1679235063
transform 1 0 15589 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_27
timestamp 1679235063
transform 1 0 15311 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_28
timestamp 1679235063
transform 1 0 19556 0 1 3336
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_29
timestamp 1679235063
transform 1 0 18631 0 1 3422
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_30
timestamp 1679235063
transform 1 0 18320 0 1 3422
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_31
timestamp 1679235063
transform 1 0 19255 0 1 3336
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_32
timestamp 1679235063
transform 1 0 18944 0 1 3336
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_33
timestamp 1679235063
transform 1 0 18198 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_34
timestamp 1679235063
transform 1 0 18476 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_35
timestamp 1679235063
transform 1 0 19374 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_36
timestamp 1679235063
transform 1 0 19100 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_37
timestamp 1679235063
transform 1 0 18788 0 1 3558
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_38
timestamp 1679235063
transform -1 0 12894 0 1 4559
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_39
timestamp 1679235063
transform 1 0 11976 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_40
timestamp 1679235063
transform 1 0 11548 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_41
timestamp 1679235063
transform 1 0 12488 0 1 4307
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_42
timestamp 1679235063
transform 1 0 13230 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_43
timestamp 1679235063
transform 1 0 12840 0 1 4313
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_44
timestamp 1679235063
transform 1 0 13386 0 -1 4805
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180857  sky130_fd_pr__via_l1m1__example_5595914180857_0
timestamp 1679235063
transform 0 1 17640 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1679235063
transform 0 -1 12402 1 0 4851
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180878  sky130_fd_pr__via_l1m1__example_5595914180878_0
timestamp 1679235063
transform -1 0 13221 0 -1 3592
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1679235063
transform 0 -1 13226 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1679235063
transform -1 0 13332 0 1 4568
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1679235063
transform 0 -1 12338 -1 0 5441
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1679235063
transform 1 0 12841 0 1 4845
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1679235063
transform 0 -1 13900 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1679235063
transform 0 -1 14836 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1679235063
transform 0 -1 14212 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1679235063
transform 0 -1 14524 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_8
timestamp 1679235063
transform 0 -1 17100 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_9
timestamp 1679235063
transform 0 -1 17412 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_10
timestamp 1679235063
transform 0 -1 20000 1 0 3638
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_11
timestamp 1679235063
transform 0 -1 19746 1 0 3638
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1679235063
transform 1 0 19591 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808291  sky130_fd_pr__via_l1m1__example_55959141808291_0
timestamp 1679235063
transform 1 0 11538 0 1 4629
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808291  sky130_fd_pr__via_l1m1__example_55959141808291_1
timestamp 1679235063
transform 1 0 11538 0 1 4771
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_0
timestamp 1679235063
transform 0 1 13498 1 0 3638
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_1
timestamp 1679235063
transform 0 1 16657 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_2
timestamp 1679235063
transform 0 1 15068 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_3
timestamp 1679235063
transform 0 1 17956 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808323  sky130_fd_pr__via_l1m1__example_55959141808323_4
timestamp 1679235063
transform 0 -1 12994 -1 0 3816
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_0
timestamp 1679235063
transform -1 0 16515 0 1 2948
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_1
timestamp 1679235063
transform 1 0 13951 0 1 3032
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808324  sky130_fd_pr__via_l1m1__example_55959141808324_2
timestamp 1679235063
transform -1 0 17944 0 1 3026
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808325  sky130_fd_pr__via_l1m1__example_55959141808325_0
timestamp 1679235063
transform 1 0 17719 0 1 4304
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1679235063
transform 1 0 11623 0 1 4155
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1679235063
transform -1 0 11651 0 1 4623
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1679235063
transform -1 0 11651 0 1 3546
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1679235063
transform -1 0 13344 0 1 4556
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1679235063
transform 1 0 13292 0 1 3020
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1679235063
transform -1 0 12600 0 1 4381
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1679235063
transform -1 0 11740 0 1 3466
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1679235063
transform -1 0 11740 0 1 4543
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1679235063
transform -1 0 13264 0 1 3020
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1679235063
transform -1 0 13264 0 1 4143
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1679235063
transform -1 0 11651 0 1 3386
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1679235063
transform 1 0 18275 0 1 3330
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_11
timestamp 1679235063
transform 0 1 13292 -1 0 3598
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_12
timestamp 1679235063
transform -1 0 18403 0 1 3020
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_13
timestamp 1679235063
transform -1 0 12600 0 1 3856
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1679235063
transform 1 0 13244 0 1 3739
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1679235063
transform 0 -1 12293 1 0 5605
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1679235063
transform 1 0 13438 0 -1 4804
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1679235063
transform 0 -1 12739 -1 0 4279
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1679235063
transform 0 -1 12904 1 0 4543
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_4
timestamp 1679235063
transform 0 -1 13091 -1 0 4279
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_5
timestamp 1679235063
transform 0 -1 13256 1 0 4543
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_6
timestamp 1679235063
transform 0 -1 13202 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_7
timestamp 1679235063
transform 0 1 13420 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_8
timestamp 1679235063
transform 0 -1 13855 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_9
timestamp 1679235063
transform 0 -1 13429 -1 0 4279
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_10
timestamp 1679235063
transform 1 0 11368 0 -1 4786
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808273  sky130_fd_pr__via_pol1__example_55959141808273_0
timestamp 1679235063
transform -1 0 12402 0 1 3252
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1679235063
transform 0 -1 13357 1 0 4105
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_0
timestamp 1679235063
transform 0 -1 18799 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_1
timestamp 1679235063
transform 0 -1 19423 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1679235063
transform 1 0 13022 0 -1 4025
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_1
timestamp 1679235063
transform 0 1 19583 1 0 4110
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808320  sky130_fd_pr__via_pol1__example_55959141808320_0
timestamp 1679235063
transform 0 -1 19265 -1 0 4354
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808321  sky130_fd_pr__via_pol1__example_55959141808321_0
timestamp 1679235063
transform 0 -1 15082 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808321  sky130_fd_pr__via_pol1__example_55959141808321_1
timestamp 1679235063
transform 0 -1 16527 -1 0 2996
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808321  sky130_fd_pr__via_pol1__example_55959141808321_2
timestamp 1679235063
transform 0 -1 17971 -1 0 3046
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808322  sky130_fd_pr__via_pol1__example_55959141808322_0
timestamp 1679235063
transform 0 1 11590 -1 0 4279
box 0 0 1 1
<< properties >>
string GDS_END 7388250
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7351164
<< end >>
