magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 13 21 1919 203
rect 25 -17 59 21
<< scnmos >>
rect 95 47 125 177
rect 179 47 209 177
rect 263 47 293 177
rect 347 47 377 177
rect 431 47 461 177
rect 515 47 545 177
rect 599 47 629 177
rect 683 47 713 177
rect 771 47 801 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1219 47 1249 177
rect 1303 47 1333 177
rect 1387 47 1417 177
rect 1471 47 1501 177
rect 1555 47 1585 177
rect 1639 47 1669 177
rect 1723 47 1753 177
rect 1807 47 1837 177
<< scpmoshvt >>
rect 95 297 125 497
rect 179 297 209 497
rect 263 297 293 497
rect 347 297 377 497
rect 431 297 461 497
rect 515 297 545 497
rect 599 297 629 497
rect 683 297 713 497
rect 871 297 901 497
rect 955 297 985 497
rect 1039 297 1069 497
rect 1123 297 1153 497
rect 1211 297 1241 497
rect 1295 297 1325 497
rect 1379 297 1409 497
rect 1463 297 1493 497
rect 1547 297 1577 497
rect 1631 297 1661 497
rect 1715 297 1745 497
rect 1799 297 1829 497
<< ndiff >>
rect 39 157 95 177
rect 39 123 51 157
rect 85 123 95 157
rect 39 89 95 123
rect 39 55 51 89
rect 85 55 95 89
rect 39 47 95 55
rect 125 129 179 177
rect 125 95 135 129
rect 169 95 179 129
rect 125 47 179 95
rect 209 89 263 177
rect 209 55 219 89
rect 253 55 263 89
rect 209 47 263 55
rect 293 129 347 177
rect 293 95 303 129
rect 337 95 347 129
rect 293 47 347 95
rect 377 89 431 177
rect 377 55 387 89
rect 421 55 431 89
rect 377 47 431 55
rect 461 129 515 177
rect 461 95 471 129
rect 505 95 515 129
rect 461 47 515 95
rect 545 89 599 177
rect 545 55 555 89
rect 589 55 599 89
rect 545 47 599 55
rect 629 129 683 177
rect 629 95 639 129
rect 673 95 683 129
rect 629 47 683 95
rect 713 89 771 177
rect 713 55 727 89
rect 761 55 771 89
rect 713 47 771 55
rect 801 129 855 177
rect 801 95 811 129
rect 845 95 855 129
rect 801 47 855 95
rect 885 89 939 177
rect 885 55 895 89
rect 929 55 939 89
rect 885 47 939 55
rect 969 129 1023 177
rect 969 95 979 129
rect 1013 95 1023 129
rect 969 47 1023 95
rect 1053 89 1109 177
rect 1053 55 1063 89
rect 1097 55 1109 89
rect 1053 47 1109 55
rect 1163 89 1219 177
rect 1163 55 1175 89
rect 1209 55 1219 89
rect 1163 47 1219 55
rect 1249 169 1303 177
rect 1249 135 1259 169
rect 1293 135 1303 169
rect 1249 47 1303 135
rect 1333 89 1387 177
rect 1333 55 1343 89
rect 1377 55 1387 89
rect 1333 47 1387 55
rect 1417 169 1471 177
rect 1417 135 1427 169
rect 1461 135 1471 169
rect 1417 47 1471 135
rect 1501 157 1555 177
rect 1501 123 1511 157
rect 1545 123 1555 157
rect 1501 89 1555 123
rect 1501 55 1511 89
rect 1545 55 1555 89
rect 1501 47 1555 55
rect 1585 169 1639 177
rect 1585 135 1595 169
rect 1629 135 1639 169
rect 1585 47 1639 135
rect 1669 89 1723 177
rect 1669 55 1679 89
rect 1713 55 1723 89
rect 1669 47 1723 55
rect 1753 169 1807 177
rect 1753 135 1763 169
rect 1797 135 1807 169
rect 1753 47 1807 135
rect 1837 89 1893 177
rect 1837 55 1847 89
rect 1881 55 1893 89
rect 1837 47 1893 55
<< pdiff >>
rect 39 448 95 497
rect 39 414 47 448
rect 81 414 95 448
rect 39 380 95 414
rect 39 346 47 380
rect 81 346 95 380
rect 39 297 95 346
rect 125 489 179 497
rect 125 455 135 489
rect 169 455 179 489
rect 125 421 179 455
rect 125 387 135 421
rect 169 387 179 421
rect 125 297 179 387
rect 209 448 263 497
rect 209 414 219 448
rect 253 414 263 448
rect 209 380 263 414
rect 209 346 219 380
rect 253 346 263 380
rect 209 297 263 346
rect 293 489 347 497
rect 293 455 303 489
rect 337 455 347 489
rect 293 421 347 455
rect 293 387 303 421
rect 337 387 347 421
rect 293 297 347 387
rect 377 448 431 497
rect 377 414 387 448
rect 421 414 431 448
rect 377 380 431 414
rect 377 346 387 380
rect 421 346 431 380
rect 377 297 431 346
rect 461 489 515 497
rect 461 455 471 489
rect 505 455 515 489
rect 461 421 515 455
rect 461 387 471 421
rect 505 387 515 421
rect 461 297 515 387
rect 545 380 599 497
rect 545 346 555 380
rect 589 346 599 380
rect 545 297 599 346
rect 629 489 683 497
rect 629 455 639 489
rect 673 455 683 489
rect 629 421 683 455
rect 629 387 639 421
rect 673 387 683 421
rect 629 297 683 387
rect 713 380 765 497
rect 713 346 723 380
rect 757 346 765 380
rect 713 297 765 346
rect 819 380 871 497
rect 819 346 827 380
rect 861 346 871 380
rect 819 297 871 346
rect 901 489 955 497
rect 901 455 911 489
rect 945 455 955 489
rect 901 421 955 455
rect 901 387 911 421
rect 945 387 955 421
rect 901 297 955 387
rect 985 380 1039 497
rect 985 346 995 380
rect 1029 346 1039 380
rect 985 297 1039 346
rect 1069 489 1123 497
rect 1069 455 1079 489
rect 1113 455 1123 489
rect 1069 421 1123 455
rect 1069 387 1079 421
rect 1113 387 1123 421
rect 1069 297 1123 387
rect 1153 448 1211 497
rect 1153 414 1163 448
rect 1197 414 1211 448
rect 1153 380 1211 414
rect 1153 346 1163 380
rect 1197 346 1211 380
rect 1153 297 1211 346
rect 1241 489 1295 497
rect 1241 455 1251 489
rect 1285 455 1295 489
rect 1241 421 1295 455
rect 1241 387 1251 421
rect 1285 387 1295 421
rect 1241 297 1295 387
rect 1325 448 1379 497
rect 1325 414 1335 448
rect 1369 414 1379 448
rect 1325 380 1379 414
rect 1325 346 1335 380
rect 1369 346 1379 380
rect 1325 297 1379 346
rect 1409 489 1463 497
rect 1409 455 1419 489
rect 1453 455 1463 489
rect 1409 421 1463 455
rect 1409 387 1419 421
rect 1453 387 1463 421
rect 1409 297 1463 387
rect 1493 448 1547 497
rect 1493 414 1503 448
rect 1537 414 1547 448
rect 1493 380 1547 414
rect 1493 346 1503 380
rect 1537 346 1547 380
rect 1493 297 1547 346
rect 1577 489 1631 497
rect 1577 455 1587 489
rect 1621 455 1631 489
rect 1577 421 1631 455
rect 1577 387 1587 421
rect 1621 387 1631 421
rect 1577 297 1631 387
rect 1661 448 1715 497
rect 1661 414 1671 448
rect 1705 414 1715 448
rect 1661 380 1715 414
rect 1661 346 1671 380
rect 1705 346 1715 380
rect 1661 297 1715 346
rect 1745 489 1799 497
rect 1745 455 1755 489
rect 1789 455 1799 489
rect 1745 421 1799 455
rect 1745 387 1755 421
rect 1789 387 1799 421
rect 1745 297 1799 387
rect 1829 448 1881 497
rect 1829 414 1839 448
rect 1873 414 1881 448
rect 1829 380 1881 414
rect 1829 346 1839 380
rect 1873 346 1881 380
rect 1829 297 1881 346
<< ndiffc >>
rect 51 123 85 157
rect 51 55 85 89
rect 135 95 169 129
rect 219 55 253 89
rect 303 95 337 129
rect 387 55 421 89
rect 471 95 505 129
rect 555 55 589 89
rect 639 95 673 129
rect 727 55 761 89
rect 811 95 845 129
rect 895 55 929 89
rect 979 95 1013 129
rect 1063 55 1097 89
rect 1175 55 1209 89
rect 1259 135 1293 169
rect 1343 55 1377 89
rect 1427 135 1461 169
rect 1511 123 1545 157
rect 1511 55 1545 89
rect 1595 135 1629 169
rect 1679 55 1713 89
rect 1763 135 1797 169
rect 1847 55 1881 89
<< pdiffc >>
rect 47 414 81 448
rect 47 346 81 380
rect 135 455 169 489
rect 135 387 169 421
rect 219 414 253 448
rect 219 346 253 380
rect 303 455 337 489
rect 303 387 337 421
rect 387 414 421 448
rect 387 346 421 380
rect 471 455 505 489
rect 471 387 505 421
rect 555 346 589 380
rect 639 455 673 489
rect 639 387 673 421
rect 723 346 757 380
rect 827 346 861 380
rect 911 455 945 489
rect 911 387 945 421
rect 995 346 1029 380
rect 1079 455 1113 489
rect 1079 387 1113 421
rect 1163 414 1197 448
rect 1163 346 1197 380
rect 1251 455 1285 489
rect 1251 387 1285 421
rect 1335 414 1369 448
rect 1335 346 1369 380
rect 1419 455 1453 489
rect 1419 387 1453 421
rect 1503 414 1537 448
rect 1503 346 1537 380
rect 1587 455 1621 489
rect 1587 387 1621 421
rect 1671 414 1705 448
rect 1671 346 1705 380
rect 1755 455 1789 489
rect 1755 387 1789 421
rect 1839 414 1873 448
rect 1839 346 1873 380
<< poly >>
rect 95 497 125 523
rect 179 497 209 523
rect 263 497 293 523
rect 347 497 377 523
rect 431 497 461 523
rect 515 497 545 523
rect 599 497 629 523
rect 683 497 713 523
rect 871 497 901 523
rect 955 497 985 523
rect 1039 497 1069 523
rect 1123 497 1153 523
rect 1211 497 1241 523
rect 1295 497 1325 523
rect 1379 497 1409 523
rect 1463 497 1493 523
rect 1547 497 1577 523
rect 1631 497 1661 523
rect 1715 497 1745 523
rect 1799 497 1829 523
rect 95 259 125 297
rect 179 259 209 297
rect 263 259 293 297
rect 347 259 377 297
rect 82 249 377 259
rect 82 215 98 249
rect 132 215 166 249
rect 200 215 234 249
rect 268 215 302 249
rect 336 215 377 249
rect 82 205 377 215
rect 95 177 125 205
rect 179 177 209 205
rect 263 177 293 205
rect 347 177 377 205
rect 431 259 461 297
rect 515 259 545 297
rect 599 259 629 297
rect 683 259 713 297
rect 871 259 901 297
rect 955 259 985 297
rect 1039 259 1069 297
rect 1123 259 1153 297
rect 431 249 713 259
rect 431 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 713 249
rect 431 205 713 215
rect 431 177 461 205
rect 515 177 545 205
rect 599 177 629 205
rect 683 177 713 205
rect 771 249 1153 259
rect 771 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 991 249
rect 1025 215 1059 249
rect 1093 215 1153 249
rect 771 205 1153 215
rect 1211 259 1241 297
rect 1295 259 1325 297
rect 1379 259 1409 297
rect 1463 259 1493 297
rect 1547 259 1577 297
rect 1631 259 1661 297
rect 1715 259 1745 297
rect 1799 259 1829 297
rect 1211 249 1501 259
rect 1211 215 1238 249
rect 1272 215 1306 249
rect 1340 215 1374 249
rect 1408 215 1442 249
rect 1476 215 1501 249
rect 1211 205 1501 215
rect 1547 249 1837 259
rect 1547 215 1589 249
rect 1623 215 1657 249
rect 1691 215 1725 249
rect 1759 215 1837 249
rect 1547 205 1837 215
rect 771 177 801 205
rect 855 177 885 205
rect 939 177 969 205
rect 1023 177 1053 205
rect 1219 177 1249 205
rect 1303 177 1333 205
rect 1387 177 1417 205
rect 1471 177 1501 205
rect 1555 177 1585 205
rect 1639 177 1669 205
rect 1723 177 1753 205
rect 1807 177 1837 205
rect 95 21 125 47
rect 179 21 209 47
rect 263 21 293 47
rect 347 21 377 47
rect 431 21 461 47
rect 515 21 545 47
rect 599 21 629 47
rect 683 21 713 47
rect 771 21 801 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1219 21 1249 47
rect 1303 21 1333 47
rect 1387 21 1417 47
rect 1471 21 1501 47
rect 1555 21 1585 47
rect 1639 21 1669 47
rect 1723 21 1753 47
rect 1807 21 1837 47
<< polycont >>
rect 98 215 132 249
rect 166 215 200 249
rect 234 215 268 249
rect 302 215 336 249
rect 447 215 481 249
rect 515 215 549 249
rect 583 215 617 249
rect 651 215 685 249
rect 787 215 821 249
rect 855 215 889 249
rect 923 215 957 249
rect 991 215 1025 249
rect 1059 215 1093 249
rect 1238 215 1272 249
rect 1306 215 1340 249
rect 1374 215 1408 249
rect 1442 215 1476 249
rect 1589 215 1623 249
rect 1657 215 1691 249
rect 1725 215 1759 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 448 81 493
rect 17 414 47 448
rect 17 380 81 414
rect 17 346 47 380
rect 119 489 185 527
rect 119 455 135 489
rect 169 455 185 489
rect 119 421 185 455
rect 119 387 135 421
rect 169 387 185 421
rect 119 379 185 387
rect 219 448 253 493
rect 219 380 253 414
rect 17 345 81 346
rect 287 489 353 527
rect 287 455 303 489
rect 337 455 353 489
rect 287 421 353 455
rect 287 387 303 421
rect 337 387 353 421
rect 287 379 353 387
rect 387 448 421 493
rect 387 380 421 414
rect 219 345 253 346
rect 455 489 1129 493
rect 455 455 471 489
rect 505 459 639 489
rect 505 455 521 459
rect 455 421 521 455
rect 623 455 639 459
rect 673 459 911 489
rect 673 455 689 459
rect 455 387 471 421
rect 505 387 521 421
rect 455 379 521 387
rect 555 380 589 423
rect 387 345 421 346
rect 623 421 689 455
rect 895 455 911 459
rect 945 459 1079 489
rect 945 455 961 459
rect 623 387 639 421
rect 673 387 689 421
rect 623 379 689 387
rect 723 380 773 423
rect 555 345 589 346
rect 757 346 773 380
rect 723 345 773 346
rect 17 297 773 345
rect 811 380 861 423
rect 811 346 827 380
rect 895 421 961 455
rect 1063 455 1079 459
rect 1113 455 1129 489
rect 895 387 911 421
rect 945 387 961 421
rect 895 379 961 387
rect 995 380 1029 423
rect 811 345 861 346
rect 1063 421 1129 455
rect 1063 387 1079 421
rect 1113 387 1129 421
rect 1063 379 1129 387
rect 1163 448 1201 493
rect 1197 414 1201 448
rect 1163 380 1201 414
rect 995 345 1029 346
rect 1197 346 1201 380
rect 1235 489 1301 527
rect 1235 455 1251 489
rect 1285 455 1301 489
rect 1235 421 1301 455
rect 1235 387 1251 421
rect 1285 387 1301 421
rect 1235 379 1301 387
rect 1335 448 1369 493
rect 1335 380 1369 414
rect 1163 345 1201 346
rect 1403 489 1469 527
rect 1403 455 1419 489
rect 1453 455 1469 489
rect 1403 421 1469 455
rect 1403 387 1419 421
rect 1453 387 1469 421
rect 1403 379 1469 387
rect 1503 448 1537 493
rect 1503 380 1537 414
rect 1335 345 1369 346
rect 1571 489 1637 527
rect 1571 455 1587 489
rect 1621 455 1637 489
rect 1571 421 1637 455
rect 1571 387 1587 421
rect 1621 387 1637 421
rect 1571 379 1637 387
rect 1671 448 1705 493
rect 1671 380 1705 414
rect 1503 345 1537 346
rect 1739 489 1805 527
rect 1739 455 1755 489
rect 1789 455 1805 489
rect 1739 421 1805 455
rect 1739 387 1755 421
rect 1789 387 1805 421
rect 1739 379 1805 387
rect 1839 448 1915 493
rect 1873 414 1915 448
rect 1839 380 1915 414
rect 1671 345 1705 346
rect 1873 346 1915 380
rect 1839 345 1915 346
rect 811 297 1915 345
rect 17 249 355 263
rect 17 215 98 249
rect 132 215 166 249
rect 200 215 234 249
rect 268 215 302 249
rect 336 215 355 249
rect 17 211 355 215
rect 389 249 723 263
rect 389 215 447 249
rect 481 215 515 249
rect 549 215 583 249
rect 617 215 651 249
rect 685 215 723 249
rect 389 211 723 215
rect 761 249 1177 263
rect 761 215 787 249
rect 821 215 855 249
rect 889 215 923 249
rect 957 215 991 249
rect 1025 215 1059 249
rect 1093 215 1177 249
rect 761 211 1177 215
rect 1211 249 1539 263
rect 1211 215 1238 249
rect 1272 215 1306 249
rect 1340 215 1374 249
rect 1408 215 1442 249
rect 1476 215 1539 249
rect 1211 211 1539 215
rect 1573 249 1818 263
rect 1573 215 1589 249
rect 1623 215 1657 249
rect 1691 215 1725 249
rect 1759 215 1818 249
rect 1573 211 1818 215
rect 1852 177 1915 297
rect 17 157 101 177
rect 17 123 51 157
rect 85 123 101 157
rect 17 89 101 123
rect 17 55 51 89
rect 85 55 101 89
rect 17 17 101 55
rect 135 169 1477 177
rect 135 135 1259 169
rect 1293 135 1427 169
rect 1461 135 1477 169
rect 135 131 1477 135
rect 1511 157 1545 177
rect 135 129 169 131
rect 303 129 337 131
rect 135 51 169 95
rect 203 89 269 97
rect 203 55 219 89
rect 253 55 269 89
rect 203 17 269 55
rect 471 129 505 131
rect 303 51 337 95
rect 371 89 437 97
rect 371 55 387 89
rect 421 55 437 89
rect 371 17 437 55
rect 639 129 673 131
rect 471 51 505 95
rect 539 89 605 97
rect 539 55 555 89
rect 589 55 605 89
rect 539 17 605 55
rect 811 129 845 131
rect 639 51 673 95
rect 707 89 777 97
rect 707 55 727 89
rect 761 55 777 89
rect 707 17 777 55
rect 979 129 1013 131
rect 811 51 845 95
rect 879 89 945 97
rect 879 55 895 89
rect 929 55 945 89
rect 879 17 945 55
rect 1579 169 1915 177
rect 1579 135 1595 169
rect 1629 135 1763 169
rect 1797 135 1915 169
rect 1579 131 1915 135
rect 1511 97 1545 123
rect 979 51 1013 95
rect 1047 89 1117 97
rect 1047 55 1063 89
rect 1097 55 1117 89
rect 1047 17 1117 55
rect 1151 89 1915 97
rect 1151 55 1175 89
rect 1209 55 1343 89
rect 1377 55 1511 89
rect 1545 55 1679 89
rect 1713 55 1847 89
rect 1881 55 1915 89
rect 1151 51 1915 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
flabel locali s 1873 425 1907 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1873 357 1907 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1873 289 1907 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1873 153 1907 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1873 221 1907 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 1781 221 1815 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1689 221 1723 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1597 221 1631 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 1505 221 1539 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1413 221 1447 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1321 221 1355 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1229 221 1263 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 1133 221 1167 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 1041 221 1075 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 949 221 983 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 857 221 891 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 765 221 799 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 669 221 703 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 577 221 611 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 485 221 519 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 393 221 427 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 301 221 335 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 209 221 243 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 117 221 151 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 25 221 59 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel metal1 s 25 -17 59 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 25 527 59 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel nwell s 25 527 59 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 25 -17 59 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 o311ai_4
rlabel metal1 s 0 -48 1932 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1932 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1932 544
string GDS_END 867278
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 851426
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.660 0.000 
<< end >>
