magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< locali >>
rect 0 1103 746 1137
rect 330 558 364 857
rect 212 485 246 551
rect 330 524 459 558
rect 557 524 591 558
rect 112 237 146 303
rect 0 -17 746 17
use pdriver  pdriver_0
timestamp 1679235063
transform 1 0 378 0 1 0
box -36 -17 404 1177
use pnand2  pnand2_0
timestamp 1679235063
transform 1 0 0 0 1 0
box -36 -17 414 1177
<< labels >>
rlabel locali s 574 541 574 541 4 Z
port 3 nsew
rlabel locali s 129 270 129 270 4 A
port 1 nsew
rlabel locali s 373 1120 373 1120 4 vdd
port 4 nsew
rlabel locali s 373 0 373 0 4 gnd
port 5 nsew
rlabel locali s 229 518 229 518 4 B
port 2 nsew
<< properties >>
string FIXED_BBOX 0 0 746 1120
string GDS_END 58022
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 56904
<< end >>
