magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 362 163 551 203
rect 1 27 551 163
rect 30 -17 64 27
rect 362 21 551 27
<< locali >>
rect 108 417 347 483
rect 481 299 535 493
rect 18 215 85 265
rect 501 152 535 299
rect 481 83 535 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 299 69 527
rect 119 265 153 377
rect 198 333 282 383
rect 383 367 439 527
rect 198 299 447 333
rect 413 265 447 299
rect 119 199 267 265
rect 413 199 459 265
rect 119 181 169 199
rect 22 147 169 181
rect 413 165 447 199
rect 22 53 84 147
rect 299 131 447 165
rect 118 17 265 113
rect 299 61 333 131
rect 367 17 443 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
rlabel locali s 108 417 347 483 6 A
port 1 nsew signal input
rlabel locali s 18 215 85 265 6 B_N
port 2 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 362 21 551 27 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 30 -17 64 27 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 27 551 163 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 362 163 551 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 481 83 535 152 6 X
port 7 nsew signal output
rlabel locali s 501 152 535 299 6 X
port 7 nsew signal output
rlabel locali s 481 299 535 493 6 X
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 999368
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 994480
<< end >>
