magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< pwell >>
rect 10 76 710 458
<< nmos >>
rect 204 102 240 432
rect 296 102 332 432
rect 388 102 424 432
rect 480 102 516 432
<< ndiff >>
rect 148 420 204 432
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 240 420 296 432
rect 240 386 251 420
rect 285 386 296 420
rect 240 352 296 386
rect 240 318 251 352
rect 285 318 296 352
rect 240 284 296 318
rect 240 250 251 284
rect 285 250 296 284
rect 240 216 296 250
rect 240 182 251 216
rect 285 182 296 216
rect 240 148 296 182
rect 240 114 251 148
rect 285 114 296 148
rect 240 102 296 114
rect 332 420 388 432
rect 332 386 343 420
rect 377 386 388 420
rect 332 352 388 386
rect 332 318 343 352
rect 377 318 388 352
rect 332 284 388 318
rect 332 250 343 284
rect 377 250 388 284
rect 332 216 388 250
rect 332 182 343 216
rect 377 182 388 216
rect 332 148 388 182
rect 332 114 343 148
rect 377 114 388 148
rect 332 102 388 114
rect 424 420 480 432
rect 424 386 435 420
rect 469 386 480 420
rect 424 352 480 386
rect 424 318 435 352
rect 469 318 480 352
rect 424 284 480 318
rect 424 250 435 284
rect 469 250 480 284
rect 424 216 480 250
rect 424 182 435 216
rect 469 182 480 216
rect 424 148 480 182
rect 424 114 435 148
rect 469 114 480 148
rect 424 102 480 114
rect 516 420 572 432
rect 516 386 527 420
rect 561 386 572 420
rect 516 352 572 386
rect 516 318 527 352
rect 561 318 572 352
rect 516 284 572 318
rect 516 250 527 284
rect 561 250 572 284
rect 516 216 572 250
rect 516 182 527 216
rect 561 182 572 216
rect 516 148 572 182
rect 516 114 527 148
rect 561 114 572 148
rect 516 102 572 114
<< ndiffc >>
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 251 386 285 420
rect 251 318 285 352
rect 251 250 285 284
rect 251 182 285 216
rect 251 114 285 148
rect 343 386 377 420
rect 343 318 377 352
rect 343 250 377 284
rect 343 182 377 216
rect 343 114 377 148
rect 435 386 469 420
rect 435 318 469 352
rect 435 250 469 284
rect 435 182 469 216
rect 435 114 469 148
rect 527 386 561 420
rect 527 318 561 352
rect 527 250 561 284
rect 527 182 561 216
rect 527 114 561 148
<< psubdiff >>
rect 36 386 94 432
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 626 386 684 432
rect 626 352 638 386
rect 672 352 684 386
rect 626 318 684 352
rect 626 284 638 318
rect 672 284 684 318
rect 626 250 684 284
rect 626 216 638 250
rect 672 216 684 250
rect 626 182 684 216
rect 626 148 638 182
rect 672 148 684 182
rect 626 102 684 148
<< psubdiffcont >>
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 638 352 672 386
rect 638 284 672 318
rect 638 216 672 250
rect 638 148 672 182
<< poly >>
rect 191 504 529 524
rect 191 470 207 504
rect 241 470 275 504
rect 309 470 343 504
rect 377 470 411 504
rect 445 470 479 504
rect 513 470 529 504
rect 191 454 529 470
rect 204 432 240 454
rect 296 432 332 454
rect 388 432 424 454
rect 480 432 516 454
rect 204 80 240 102
rect 296 80 332 102
rect 388 80 424 102
rect 480 80 516 102
rect 191 64 529 80
rect 191 30 207 64
rect 241 30 275 64
rect 309 30 343 64
rect 377 30 411 64
rect 445 30 479 64
rect 513 30 529 64
rect 191 10 529 30
<< polycont >>
rect 207 470 241 504
rect 275 470 309 504
rect 343 470 377 504
rect 411 470 445 504
rect 479 470 513 504
rect 207 30 241 64
rect 275 30 309 64
rect 343 30 377 64
rect 411 30 445 64
rect 479 30 513 64
<< locali >>
rect 191 470 199 504
rect 241 470 271 504
rect 309 470 343 504
rect 377 470 411 504
rect 449 470 479 504
rect 521 470 529 504
rect 159 420 193 436
rect 48 392 82 402
rect 48 320 82 352
rect 48 250 82 284
rect 48 182 82 214
rect 48 132 82 142
rect 159 352 193 358
rect 159 284 193 286
rect 159 248 193 250
rect 159 176 193 182
rect 159 98 193 114
rect 251 420 285 436
rect 251 352 285 358
rect 251 284 285 286
rect 251 248 285 250
rect 251 176 285 182
rect 251 98 285 114
rect 343 420 377 436
rect 343 352 377 358
rect 343 284 377 286
rect 343 248 377 250
rect 343 176 377 182
rect 343 98 377 114
rect 435 420 469 436
rect 435 352 469 358
rect 435 284 469 286
rect 435 248 469 250
rect 435 176 469 182
rect 435 98 469 114
rect 527 420 561 436
rect 527 352 561 358
rect 527 284 561 286
rect 527 248 561 250
rect 527 176 561 182
rect 638 392 672 402
rect 638 320 672 352
rect 638 250 672 284
rect 638 182 672 214
rect 638 132 672 142
rect 527 98 561 114
rect 191 30 199 64
rect 241 30 271 64
rect 309 30 343 64
rect 377 30 411 64
rect 449 30 479 64
rect 521 30 529 64
<< viali >>
rect 199 470 207 504
rect 207 470 233 504
rect 271 470 275 504
rect 275 470 305 504
rect 343 470 377 504
rect 415 470 445 504
rect 445 470 449 504
rect 487 470 513 504
rect 513 470 521 504
rect 48 386 82 392
rect 48 358 82 386
rect 48 318 82 320
rect 48 286 82 318
rect 48 216 82 248
rect 48 214 82 216
rect 48 148 82 176
rect 48 142 82 148
rect 159 386 193 392
rect 159 358 193 386
rect 159 318 193 320
rect 159 286 193 318
rect 159 216 193 248
rect 159 214 193 216
rect 159 148 193 176
rect 159 142 193 148
rect 251 386 285 392
rect 251 358 285 386
rect 251 318 285 320
rect 251 286 285 318
rect 251 216 285 248
rect 251 214 285 216
rect 251 148 285 176
rect 251 142 285 148
rect 343 386 377 392
rect 343 358 377 386
rect 343 318 377 320
rect 343 286 377 318
rect 343 216 377 248
rect 343 214 377 216
rect 343 148 377 176
rect 343 142 377 148
rect 435 386 469 392
rect 435 358 469 386
rect 435 318 469 320
rect 435 286 469 318
rect 435 216 469 248
rect 435 214 469 216
rect 435 148 469 176
rect 435 142 469 148
rect 527 386 561 392
rect 527 358 561 386
rect 527 318 561 320
rect 527 286 561 318
rect 527 216 561 248
rect 527 214 561 216
rect 527 148 561 176
rect 527 142 561 148
rect 638 386 672 392
rect 638 358 672 386
rect 638 318 672 320
rect 638 286 672 318
rect 638 216 672 248
rect 638 214 672 216
rect 638 148 672 176
rect 638 142 672 148
rect 199 30 207 64
rect 207 30 233 64
rect 271 30 275 64
rect 275 30 305 64
rect 343 30 377 64
rect 415 30 445 64
rect 445 30 449 64
rect 487 30 513 64
rect 513 30 521 64
<< metal1 >>
rect 187 504 533 524
rect 187 470 199 504
rect 233 470 271 504
rect 305 470 343 504
rect 377 470 415 504
rect 449 470 487 504
rect 521 470 533 504
rect 187 458 533 470
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 150 392 202 420
rect 150 358 159 392
rect 193 358 202 392
rect 150 320 202 358
rect 150 286 159 320
rect 193 286 202 320
rect 150 248 202 286
rect 150 236 159 248
rect 193 236 202 248
rect 150 176 202 184
rect 150 172 159 176
rect 193 172 202 176
rect 150 114 202 120
rect 242 414 294 420
rect 242 358 251 362
rect 285 358 294 362
rect 242 350 294 358
rect 242 286 251 298
rect 285 286 294 298
rect 242 248 294 286
rect 242 214 251 248
rect 285 214 294 248
rect 242 176 294 214
rect 242 142 251 176
rect 285 142 294 176
rect 242 114 294 142
rect 334 392 386 420
rect 334 358 343 392
rect 377 358 386 392
rect 334 320 386 358
rect 334 286 343 320
rect 377 286 386 320
rect 334 248 386 286
rect 334 236 343 248
rect 377 236 386 248
rect 334 176 386 184
rect 334 172 343 176
rect 377 172 386 176
rect 334 114 386 120
rect 426 414 478 420
rect 426 358 435 362
rect 469 358 478 362
rect 426 350 478 358
rect 426 286 435 298
rect 469 286 478 298
rect 426 248 478 286
rect 426 214 435 248
rect 469 214 478 248
rect 426 176 478 214
rect 426 142 435 176
rect 469 142 478 176
rect 426 114 478 142
rect 518 392 570 420
rect 518 358 527 392
rect 561 358 570 392
rect 518 320 570 358
rect 518 286 527 320
rect 561 286 570 320
rect 518 248 570 286
rect 518 236 527 248
rect 561 236 570 248
rect 518 176 570 184
rect 518 172 527 176
rect 561 172 570 176
rect 518 114 570 120
rect 626 392 684 420
rect 626 358 638 392
rect 672 358 684 392
rect 626 320 684 358
rect 626 286 638 320
rect 672 286 684 320
rect 626 248 684 286
rect 626 214 638 248
rect 672 214 684 248
rect 626 176 684 214
rect 626 142 638 176
rect 672 142 684 176
rect 626 114 684 142
rect 187 64 533 76
rect 187 30 199 64
rect 233 30 271 64
rect 305 30 343 64
rect 377 30 415 64
rect 449 30 487 64
rect 521 30 533 64
rect 187 10 533 30
<< via1 >>
rect 150 214 159 236
rect 159 214 193 236
rect 193 214 202 236
rect 150 184 202 214
rect 150 142 159 172
rect 159 142 193 172
rect 193 142 202 172
rect 150 120 202 142
rect 242 392 294 414
rect 242 362 251 392
rect 251 362 285 392
rect 285 362 294 392
rect 242 320 294 350
rect 242 298 251 320
rect 251 298 285 320
rect 285 298 294 320
rect 334 214 343 236
rect 343 214 377 236
rect 377 214 386 236
rect 334 184 386 214
rect 334 142 343 172
rect 343 142 377 172
rect 377 142 386 172
rect 334 120 386 142
rect 426 392 478 414
rect 426 362 435 392
rect 435 362 469 392
rect 469 362 478 392
rect 426 320 478 350
rect 426 298 435 320
rect 435 298 469 320
rect 469 298 478 320
rect 518 214 527 236
rect 527 214 561 236
rect 561 214 570 236
rect 518 184 570 214
rect 518 142 527 172
rect 527 142 561 172
rect 561 142 570 172
rect 518 120 570 142
<< metal2 >>
rect 10 414 710 420
rect 10 362 242 414
rect 294 362 426 414
rect 478 362 710 414
rect 10 350 710 362
rect 10 298 242 350
rect 294 298 426 350
rect 478 298 710 350
rect 10 292 710 298
rect 10 236 710 242
rect 10 184 150 236
rect 202 184 334 236
rect 386 184 518 236
rect 570 184 710 236
rect 10 172 710 184
rect 10 120 150 172
rect 202 120 334 172
rect 386 120 518 172
rect 570 120 710 172
rect 10 114 710 120
<< labels >>
flabel metal2 s 10 292 30 420 7 FreeSans 300 180 0 0 DRAIN
port 2 nsew
flabel metal2 s 10 114 30 242 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal1 s 187 10 533 76 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 187 458 533 524 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 626 114 684 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
flabel metal1 s 36 114 94 130 3 FreeSans 300 90 0 0 SUBSTRATE
port 5 nsew
<< properties >>
string GDS_END 5016034
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5005638
<< end >>
