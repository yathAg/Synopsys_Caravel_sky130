magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 99 157 509 203
rect 1 21 721 157
rect 29 -17 63 21
<< scnmos >>
rect 80 47 110 131
rect 175 47 225 177
rect 383 47 433 177
rect 498 47 528 131
rect 598 47 628 131
<< scpmoshvt >>
rect 80 297 110 497
rect 175 333 225 497
rect 383 333 433 497
rect 498 297 528 497
rect 598 297 628 497
<< ndiff >>
rect 125 131 175 177
rect 27 111 80 131
rect 27 77 35 111
rect 69 77 80 111
rect 27 47 80 77
rect 110 94 175 131
rect 110 60 131 94
rect 165 60 175 94
rect 110 47 175 60
rect 225 120 277 177
rect 225 86 235 120
rect 269 86 277 120
rect 225 47 277 86
rect 331 99 383 177
rect 331 65 339 99
rect 373 65 383 99
rect 331 47 383 65
rect 433 131 483 177
rect 433 93 498 131
rect 433 59 443 93
rect 477 59 498 93
rect 433 47 498 59
rect 528 107 598 131
rect 528 73 554 107
rect 588 73 598 107
rect 528 47 598 73
rect 628 94 695 131
rect 628 60 653 94
rect 687 60 695 94
rect 628 47 695 60
<< pdiff >>
rect 27 475 80 497
rect 27 441 35 475
rect 69 441 80 475
rect 27 407 80 441
rect 27 373 35 407
rect 69 373 80 407
rect 27 297 80 373
rect 110 485 175 497
rect 110 451 131 485
rect 165 451 175 485
rect 110 333 175 451
rect 225 477 277 497
rect 225 443 235 477
rect 269 443 277 477
rect 225 379 277 443
rect 225 345 235 379
rect 269 345 277 379
rect 225 333 277 345
rect 331 477 383 497
rect 331 443 339 477
rect 373 443 383 477
rect 331 379 383 443
rect 331 345 339 379
rect 373 345 383 379
rect 331 333 383 345
rect 433 485 498 497
rect 433 451 443 485
rect 477 451 498 485
rect 433 417 498 451
rect 433 383 443 417
rect 477 383 498 417
rect 433 333 498 383
rect 110 297 160 333
rect 448 297 498 333
rect 528 476 598 497
rect 528 442 554 476
rect 588 442 598 476
rect 528 375 598 442
rect 528 341 554 375
rect 588 341 598 375
rect 528 297 598 341
rect 628 485 695 497
rect 628 451 653 485
rect 687 451 695 485
rect 628 388 695 451
rect 628 354 653 388
rect 687 354 695 388
rect 628 297 695 354
<< ndiffc >>
rect 35 77 69 111
rect 131 60 165 94
rect 235 86 269 120
rect 339 65 373 99
rect 443 59 477 93
rect 554 73 588 107
rect 653 60 687 94
<< pdiffc >>
rect 35 441 69 475
rect 35 373 69 407
rect 131 451 165 485
rect 235 443 269 477
rect 235 345 269 379
rect 339 443 373 477
rect 339 345 373 379
rect 443 451 477 485
rect 443 383 477 417
rect 554 442 588 476
rect 554 341 588 375
rect 653 451 687 485
rect 653 354 687 388
<< poly >>
rect 80 497 110 523
rect 175 497 225 523
rect 383 497 433 523
rect 498 497 528 523
rect 598 497 628 523
rect 80 265 110 297
rect 175 265 225 333
rect 383 265 433 333
rect 498 268 528 297
rect 598 268 628 297
rect 498 265 628 268
rect 44 249 110 265
rect 44 215 54 249
rect 88 215 110 249
rect 44 194 110 215
rect 163 249 225 265
rect 163 215 173 249
rect 207 215 225 249
rect 163 199 225 215
rect 275 249 433 265
rect 275 215 285 249
rect 319 215 389 249
rect 423 215 433 249
rect 275 199 433 215
rect 475 249 628 265
rect 475 215 485 249
rect 519 215 628 249
rect 475 199 628 215
rect 80 131 110 194
rect 175 177 225 199
rect 383 177 433 199
rect 498 197 628 199
rect 498 131 528 197
rect 598 131 628 197
rect 80 21 110 47
rect 175 21 225 47
rect 383 21 433 47
rect 498 21 528 47
rect 598 21 628 47
<< polycont >>
rect 54 215 88 249
rect 173 215 207 249
rect 285 215 319 249
rect 389 215 423 249
rect 485 215 519 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 19 475 69 493
rect 19 441 35 475
rect 19 407 69 441
rect 115 485 181 527
rect 115 451 131 485
rect 165 451 181 485
rect 115 425 181 451
rect 235 477 288 493
rect 269 443 288 477
rect 19 373 35 407
rect 69 373 167 391
rect 19 357 167 373
rect 133 350 167 357
rect 235 379 288 443
rect 17 249 99 323
rect 17 215 54 249
rect 88 215 99 249
rect 17 199 99 215
rect 133 265 201 350
rect 269 345 288 379
rect 235 285 288 345
rect 339 477 389 493
rect 373 443 389 477
rect 339 379 389 443
rect 427 485 493 527
rect 427 451 443 485
rect 477 451 493 485
rect 427 417 493 451
rect 427 383 443 417
rect 477 383 493 417
rect 554 476 619 492
rect 588 442 619 476
rect 373 349 389 379
rect 554 375 619 442
rect 373 345 519 349
rect 339 300 519 345
rect 588 341 619 375
rect 554 325 619 341
rect 653 485 719 527
rect 687 451 719 485
rect 653 388 719 451
rect 687 354 719 388
rect 653 327 719 354
rect 241 265 288 285
rect 133 249 207 265
rect 133 215 173 249
rect 133 199 207 215
rect 241 249 433 265
rect 241 215 285 249
rect 319 215 389 249
rect 423 215 433 249
rect 241 199 433 215
rect 467 249 519 300
rect 467 215 485 249
rect 133 162 168 199
rect 19 128 168 162
rect 241 156 285 199
rect 467 161 519 215
rect 19 111 69 128
rect 19 77 35 111
rect 219 120 285 156
rect 19 61 69 77
rect 115 60 131 94
rect 165 60 181 94
rect 115 17 181 60
rect 219 86 235 120
rect 269 86 285 120
rect 219 51 285 86
rect 323 127 519 161
rect 573 255 619 325
rect 573 153 719 255
rect 323 99 389 127
rect 573 123 619 153
rect 323 65 339 99
rect 373 65 389 99
rect 554 107 619 123
rect 323 51 389 65
rect 427 59 443 93
rect 477 59 493 93
rect 427 17 493 59
rect 588 73 619 107
rect 554 57 619 73
rect 653 94 719 110
rect 687 60 719 94
rect 653 17 719 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 585 221 619 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 585 85 619 119 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 585 425 619 459 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 677 153 711 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 585 153 619 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 585 357 619 391 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 677 221 711 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 clkdlybuf4s25_2
rlabel metal1 s 0 -48 736 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3290926
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3284314
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 18.400 13.600 
<< end >>
