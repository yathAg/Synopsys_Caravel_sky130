magic
tech sky130A
magscale 1 2
timestamp 1679235063
use sky130_fd_io__gpiov2_amux_decoder  sky130_fd_io__gpiov2_amux_decoder_0
timestamp 1679235063
transform 1 0 31774 0 1 -5388
box 362 211 8121 2886
use sky130_fd_io__gpiov2_amux_drvr  sky130_fd_io__gpiov2_amux_drvr_0
timestamp 1679235063
transform 1 0 9862 0 1 6253
box 16319 -13467 28102 -4405
use sky130_fd_io__gpiov2_amux_ls  sky130_fd_io__gpiov2_amux_ls_0
timestamp 1679235063
transform 1 0 25054 0 1 -16031
box 1038 445 16816 16947
<< properties >>
string GDS_END 8666320
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8597136
<< end >>
