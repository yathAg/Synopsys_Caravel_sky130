magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< locali >>
rect 383 961 667 980
rect 383 855 400 961
rect 650 855 667 961
rect 383 843 667 855
rect 383 125 667 137
rect 383 19 400 125
rect 650 19 667 125
rect 383 0 667 19
<< viali >>
rect 400 855 650 961
rect 400 19 650 125
<< obsli1 >>
rect 190 817 256 883
rect 794 817 860 883
rect 190 795 230 817
rect 820 795 860 817
rect 41 759 230 795
rect 41 725 60 759
rect 94 725 230 759
rect 41 687 230 725
rect 41 653 60 687
rect 94 653 230 687
rect 41 615 230 653
rect 41 581 60 615
rect 94 581 230 615
rect 41 543 230 581
rect 41 509 60 543
rect 94 509 230 543
rect 41 471 230 509
rect 41 437 60 471
rect 94 437 230 471
rect 41 399 230 437
rect 41 365 60 399
rect 94 365 230 399
rect 41 327 230 365
rect 41 293 60 327
rect 94 293 230 327
rect 41 255 230 293
rect 41 221 60 255
rect 94 221 230 255
rect 41 185 230 221
rect 352 185 386 795
rect 508 185 542 795
rect 664 185 698 795
rect 820 759 1009 795
rect 820 725 956 759
rect 990 725 1009 759
rect 820 687 1009 725
rect 820 653 956 687
rect 990 653 1009 687
rect 820 615 1009 653
rect 820 581 956 615
rect 990 581 1009 615
rect 820 543 1009 581
rect 820 509 956 543
rect 990 509 1009 543
rect 820 471 1009 509
rect 820 437 956 471
rect 990 437 1009 471
rect 820 399 1009 437
rect 820 365 956 399
rect 990 365 1009 399
rect 820 327 1009 365
rect 820 293 956 327
rect 990 293 1009 327
rect 820 255 1009 293
rect 820 221 956 255
rect 990 221 1009 255
rect 820 185 1009 221
rect 190 163 230 185
rect 820 163 860 185
rect 190 97 256 163
rect 794 97 860 163
<< obsli1c >>
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 956 725 990 759
rect 956 653 990 687
rect 956 581 990 615
rect 956 509 990 543
rect 956 437 990 471
rect 956 365 990 399
rect 956 293 990 327
rect 956 221 990 255
<< metal1 >>
rect 380 961 670 980
rect 380 855 400 961
rect 650 855 670 961
rect 380 843 670 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 950 759 1009 771
rect 950 725 956 759
rect 990 725 1009 759
rect 950 687 1009 725
rect 950 653 956 687
rect 990 653 1009 687
rect 950 615 1009 653
rect 950 581 956 615
rect 990 581 1009 615
rect 950 543 1009 581
rect 950 509 956 543
rect 990 509 1009 543
rect 950 471 1009 509
rect 950 437 956 471
rect 990 437 1009 471
rect 950 399 1009 437
rect 950 365 956 399
rect 990 365 1009 399
rect 950 327 1009 365
rect 950 293 956 327
rect 990 293 1009 327
rect 950 255 1009 293
rect 950 221 956 255
rect 990 221 1009 255
rect 950 209 1009 221
rect 380 125 670 137
rect 380 19 400 125
rect 650 19 670 125
rect 380 0 670 19
<< obsm1 >>
rect 343 209 395 771
rect 499 209 551 771
rect 655 209 707 771
<< metal2 >>
rect 14 515 1036 771
rect 14 209 1036 465
<< labels >>
rlabel metal2 s 14 515 1036 771 6 DRAIN
port 1 nsew
rlabel viali s 400 855 650 961 6 GATE
port 2 nsew
rlabel viali s 400 19 650 125 6 GATE
port 2 nsew
rlabel locali s 383 843 667 980 6 GATE
port 2 nsew
rlabel locali s 383 0 667 137 6 GATE
port 2 nsew
rlabel metal1 s 380 843 670 980 6 GATE
port 2 nsew
rlabel metal1 s 380 0 670 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 1036 465 6 SOURCE
port 3 nsew
rlabel metal1 s 41 209 100 771 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 950 209 1009 771 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 1036 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7645460
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7628736
string device primitive
<< end >>
