magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< dnwell >>
rect -1298 -1522 1448 7522
<< nwell >>
rect -898 6600 1048 7122
rect -898 6026 -500 6600
rect 650 6026 1048 6600
rect -898 -26 -526 6026
rect 676 -26 1048 6026
rect -898 -600 -500 -26
rect 650 -600 1048 -26
rect -898 -1122 1048 -600
<< pwell >>
rect -1606 7696 1756 7830
rect -1606 -1696 -1472 7696
rect -526 -26 -274 6026
tri -26 5996 4 6026 se
rect 4 5996 146 6026
tri 146 5996 176 6026 sw
rect -26 4 176 5996
tri -26 -26 4 4 ne
rect 4 -26 146 4
tri 146 -26 176 4 nw
rect 424 -26 676 6026
rect 1622 -1696 1756 7696
rect -1606 -1830 1756 -1696
<< obsactive >>
rect -1730 -1954 1880 7954
<< locali >>
rect -1580 7780 1730 7804
rect -1580 7746 -1454 7780
rect -1420 7746 -1382 7780
rect -1348 7746 -1310 7780
rect -1276 7746 -1238 7780
rect -1204 7746 -1166 7780
rect -1132 7746 -1094 7780
rect -1060 7746 -1022 7780
rect -988 7746 -950 7780
rect -916 7746 -878 7780
rect -844 7746 -806 7780
rect -772 7746 -734 7780
rect -700 7746 -662 7780
rect -628 7746 -590 7780
rect -556 7746 -518 7780
rect -484 7746 -446 7780
rect -412 7746 -374 7780
rect -340 7746 -302 7780
rect -268 7746 -230 7780
rect -196 7746 -158 7780
rect -124 7746 -86 7780
rect -52 7746 -14 7780
rect 20 7746 58 7780
rect 92 7746 130 7780
rect 164 7746 202 7780
rect 236 7746 274 7780
rect 308 7746 346 7780
rect 380 7746 418 7780
rect 452 7746 490 7780
rect 524 7746 562 7780
rect 596 7746 634 7780
rect 668 7746 706 7780
rect 740 7746 778 7780
rect 812 7746 850 7780
rect 884 7746 922 7780
rect 956 7746 994 7780
rect 1028 7746 1066 7780
rect 1100 7746 1138 7780
rect 1172 7746 1210 7780
rect 1244 7746 1282 7780
rect 1316 7746 1354 7780
rect 1388 7746 1426 7780
rect 1460 7746 1498 7780
rect 1532 7746 1570 7780
rect 1604 7746 1730 7780
rect -1580 7722 1730 7746
rect -1580 7661 -1498 7722
rect -1580 7627 -1556 7661
rect -1522 7627 -1498 7661
rect -1580 7589 -1498 7627
rect -1580 7555 -1556 7589
rect -1522 7555 -1498 7589
rect -1580 7517 -1498 7555
rect -1580 7483 -1556 7517
rect -1522 7483 -1498 7517
rect -1580 7445 -1498 7483
rect -1580 7411 -1556 7445
rect -1522 7411 -1498 7445
rect -1580 7373 -1498 7411
rect -1580 7339 -1556 7373
rect -1522 7339 -1498 7373
rect -1580 7301 -1498 7339
rect -1580 7267 -1556 7301
rect -1522 7267 -1498 7301
rect -1580 7229 -1498 7267
rect -1580 7195 -1556 7229
rect -1522 7195 -1498 7229
rect -1580 7157 -1498 7195
rect -1580 7123 -1556 7157
rect -1522 7123 -1498 7157
rect -1580 7085 -1498 7123
rect -1580 7051 -1556 7085
rect -1522 7051 -1498 7085
rect -1580 7013 -1498 7051
rect 1648 7661 1730 7722
rect 1648 7627 1672 7661
rect 1706 7627 1730 7661
rect 1648 7589 1730 7627
rect 1648 7555 1672 7589
rect 1706 7555 1730 7589
rect 1648 7517 1730 7555
rect 1648 7483 1672 7517
rect 1706 7483 1730 7517
rect 1648 7445 1730 7483
rect 1648 7411 1672 7445
rect 1706 7411 1730 7445
rect 1648 7373 1730 7411
rect 1648 7339 1672 7373
rect 1706 7339 1730 7373
rect 1648 7301 1730 7339
rect 1648 7267 1672 7301
rect 1706 7267 1730 7301
rect 1648 7229 1730 7267
rect 1648 7195 1672 7229
rect 1706 7195 1730 7229
rect 1648 7157 1730 7195
rect 1648 7123 1672 7157
rect 1706 7123 1730 7157
rect 1648 7085 1730 7123
rect 1648 7051 1672 7085
rect 1706 7051 1730 7085
rect -1580 6979 -1556 7013
rect -1522 6979 -1498 7013
rect -1580 6941 -1498 6979
rect -1580 6907 -1556 6941
rect -1522 6907 -1498 6941
rect -1580 6869 -1498 6907
rect -1580 6835 -1556 6869
rect -1522 6835 -1498 6869
rect -1580 6797 -1498 6835
rect -1580 6763 -1556 6797
rect -1522 6763 -1498 6797
rect -1580 6725 -1498 6763
rect -1580 6691 -1556 6725
rect -1522 6691 -1498 6725
rect -1580 6653 -1498 6691
rect -1580 6619 -1556 6653
rect -1522 6619 -1498 6653
rect -1580 6581 -1498 6619
rect -1580 6547 -1556 6581
rect -1522 6547 -1498 6581
rect -1580 6509 -1498 6547
rect -1580 6475 -1556 6509
rect -1522 6475 -1498 6509
rect -1580 6437 -1498 6475
rect -1580 6403 -1556 6437
rect -1522 6403 -1498 6437
rect -1580 6365 -1498 6403
rect -1580 6331 -1556 6365
rect -1522 6331 -1498 6365
rect -1580 6293 -1498 6331
rect -1580 6259 -1556 6293
rect -1522 6259 -1498 6293
rect -1580 6221 -1498 6259
rect -1580 6187 -1556 6221
rect -1522 6187 -1498 6221
rect -1580 6149 -1498 6187
rect -1580 6115 -1556 6149
rect -1522 6115 -1498 6149
rect -1580 6077 -1498 6115
rect -1580 6043 -1556 6077
rect -1522 6043 -1498 6077
rect -1580 6005 -1498 6043
rect -1580 5971 -1556 6005
rect -1522 5971 -1498 6005
rect -1580 5933 -1498 5971
rect -1580 5899 -1556 5933
rect -1522 5899 -1498 5933
rect -1580 5861 -1498 5899
rect -1580 5827 -1556 5861
rect -1522 5827 -1498 5861
rect -1580 5789 -1498 5827
rect -1580 5755 -1556 5789
rect -1522 5755 -1498 5789
rect -1580 5717 -1498 5755
rect -1580 5683 -1556 5717
rect -1522 5683 -1498 5717
rect -1580 5645 -1498 5683
rect -1580 5611 -1556 5645
rect -1522 5611 -1498 5645
rect -1580 5573 -1498 5611
rect -1580 5539 -1556 5573
rect -1522 5539 -1498 5573
rect -1580 5501 -1498 5539
rect -1580 5467 -1556 5501
rect -1522 5467 -1498 5501
rect -1580 5429 -1498 5467
rect -1580 5395 -1556 5429
rect -1522 5395 -1498 5429
rect -1580 5357 -1498 5395
rect -1580 5323 -1556 5357
rect -1522 5323 -1498 5357
rect -1580 5285 -1498 5323
rect -1580 5251 -1556 5285
rect -1522 5251 -1498 5285
rect -1580 5213 -1498 5251
rect -1580 5179 -1556 5213
rect -1522 5179 -1498 5213
rect -1580 5141 -1498 5179
rect -1580 5107 -1556 5141
rect -1522 5107 -1498 5141
rect -1580 5069 -1498 5107
rect -1580 5035 -1556 5069
rect -1522 5035 -1498 5069
rect -1580 4997 -1498 5035
rect -1580 4963 -1556 4997
rect -1522 4963 -1498 4997
rect -1580 4925 -1498 4963
rect -1580 4891 -1556 4925
rect -1522 4891 -1498 4925
rect -1580 4853 -1498 4891
rect -1580 4819 -1556 4853
rect -1522 4819 -1498 4853
rect -1580 4781 -1498 4819
rect -1580 4747 -1556 4781
rect -1522 4747 -1498 4781
rect -1580 4709 -1498 4747
rect -1580 4675 -1556 4709
rect -1522 4675 -1498 4709
rect -1580 4637 -1498 4675
rect -1580 4603 -1556 4637
rect -1522 4603 -1498 4637
rect -1580 4565 -1498 4603
rect -1580 4531 -1556 4565
rect -1522 4531 -1498 4565
rect -1580 4493 -1498 4531
rect -1580 4459 -1556 4493
rect -1522 4459 -1498 4493
rect -1580 4421 -1498 4459
rect -1580 4387 -1556 4421
rect -1522 4387 -1498 4421
rect -1580 4349 -1498 4387
rect -1580 4315 -1556 4349
rect -1522 4315 -1498 4349
rect -1580 4277 -1498 4315
rect -1580 4243 -1556 4277
rect -1522 4243 -1498 4277
rect -1580 4205 -1498 4243
rect -1580 4171 -1556 4205
rect -1522 4171 -1498 4205
rect -1580 4133 -1498 4171
rect -1580 4099 -1556 4133
rect -1522 4099 -1498 4133
rect -1580 4061 -1498 4099
rect -1580 4027 -1556 4061
rect -1522 4027 -1498 4061
rect -1580 3989 -1498 4027
rect -1580 3955 -1556 3989
rect -1522 3955 -1498 3989
rect -1580 3917 -1498 3955
rect -1580 3883 -1556 3917
rect -1522 3883 -1498 3917
rect -1580 3845 -1498 3883
rect -1580 3811 -1556 3845
rect -1522 3811 -1498 3845
rect -1580 3773 -1498 3811
rect -1580 3739 -1556 3773
rect -1522 3739 -1498 3773
rect -1580 3701 -1498 3739
rect -1580 3667 -1556 3701
rect -1522 3667 -1498 3701
rect -1580 3629 -1498 3667
rect -1580 3595 -1556 3629
rect -1522 3595 -1498 3629
rect -1580 3557 -1498 3595
rect -1580 3523 -1556 3557
rect -1522 3523 -1498 3557
rect -1580 3485 -1498 3523
rect -1580 3451 -1556 3485
rect -1522 3451 -1498 3485
rect -1580 3413 -1498 3451
rect -1580 3379 -1556 3413
rect -1522 3379 -1498 3413
rect -1580 3341 -1498 3379
rect -1580 3307 -1556 3341
rect -1522 3307 -1498 3341
rect -1580 3269 -1498 3307
rect -1580 3235 -1556 3269
rect -1522 3235 -1498 3269
rect -1580 3197 -1498 3235
rect -1580 3163 -1556 3197
rect -1522 3163 -1498 3197
rect -1580 3125 -1498 3163
rect -1580 3091 -1556 3125
rect -1522 3091 -1498 3125
rect -1580 3053 -1498 3091
rect -1580 3019 -1556 3053
rect -1522 3019 -1498 3053
rect -1580 2981 -1498 3019
rect -1580 2947 -1556 2981
rect -1522 2947 -1498 2981
rect -1580 2909 -1498 2947
rect -1580 2875 -1556 2909
rect -1522 2875 -1498 2909
rect -1580 2837 -1498 2875
rect -1580 2803 -1556 2837
rect -1522 2803 -1498 2837
rect -1580 2765 -1498 2803
rect -1580 2731 -1556 2765
rect -1522 2731 -1498 2765
rect -1580 2693 -1498 2731
rect -1580 2659 -1556 2693
rect -1522 2659 -1498 2693
rect -1580 2621 -1498 2659
rect -1580 2587 -1556 2621
rect -1522 2587 -1498 2621
rect -1580 2549 -1498 2587
rect -1580 2515 -1556 2549
rect -1522 2515 -1498 2549
rect -1580 2477 -1498 2515
rect -1580 2443 -1556 2477
rect -1522 2443 -1498 2477
rect -1580 2405 -1498 2443
rect -1580 2371 -1556 2405
rect -1522 2371 -1498 2405
rect -1580 2333 -1498 2371
rect -1580 2299 -1556 2333
rect -1522 2299 -1498 2333
rect -1580 2261 -1498 2299
rect -1580 2227 -1556 2261
rect -1522 2227 -1498 2261
rect -1580 2189 -1498 2227
rect -1580 2155 -1556 2189
rect -1522 2155 -1498 2189
rect -1580 2117 -1498 2155
rect -1580 2083 -1556 2117
rect -1522 2083 -1498 2117
rect -1580 2045 -1498 2083
rect -1580 2011 -1556 2045
rect -1522 2011 -1498 2045
rect -1580 1973 -1498 2011
rect -1580 1939 -1556 1973
rect -1522 1939 -1498 1973
rect -1580 1901 -1498 1939
rect -1580 1867 -1556 1901
rect -1522 1867 -1498 1901
rect -1580 1829 -1498 1867
rect -1580 1795 -1556 1829
rect -1522 1795 -1498 1829
rect -1580 1757 -1498 1795
rect -1580 1723 -1556 1757
rect -1522 1723 -1498 1757
rect -1580 1685 -1498 1723
rect -1580 1651 -1556 1685
rect -1522 1651 -1498 1685
rect -1580 1613 -1498 1651
rect -1580 1579 -1556 1613
rect -1522 1579 -1498 1613
rect -1580 1541 -1498 1579
rect -1580 1507 -1556 1541
rect -1522 1507 -1498 1541
rect -1580 1469 -1498 1507
rect -1580 1435 -1556 1469
rect -1522 1435 -1498 1469
rect -1580 1397 -1498 1435
rect -1580 1363 -1556 1397
rect -1522 1363 -1498 1397
rect -1580 1325 -1498 1363
rect -1580 1291 -1556 1325
rect -1522 1291 -1498 1325
rect -1580 1253 -1498 1291
rect -1580 1219 -1556 1253
rect -1522 1219 -1498 1253
rect -1580 1181 -1498 1219
rect -1580 1147 -1556 1181
rect -1522 1147 -1498 1181
rect -1580 1109 -1498 1147
rect -1580 1075 -1556 1109
rect -1522 1075 -1498 1109
rect -1580 1037 -1498 1075
rect -1580 1003 -1556 1037
rect -1522 1003 -1498 1037
rect -1580 965 -1498 1003
rect -1580 931 -1556 965
rect -1522 931 -1498 965
rect -1580 893 -1498 931
rect -1580 859 -1556 893
rect -1522 859 -1498 893
rect -1580 821 -1498 859
rect -1580 787 -1556 821
rect -1522 787 -1498 821
rect -1580 749 -1498 787
rect -1580 715 -1556 749
rect -1522 715 -1498 749
rect -1580 677 -1498 715
rect -1580 643 -1556 677
rect -1522 643 -1498 677
rect -1580 605 -1498 643
rect -1580 571 -1556 605
rect -1522 571 -1498 605
rect -1580 533 -1498 571
rect -1580 499 -1556 533
rect -1522 499 -1498 533
rect -1580 461 -1498 499
rect -1580 427 -1556 461
rect -1522 427 -1498 461
rect -1580 389 -1498 427
rect -1580 355 -1556 389
rect -1522 355 -1498 389
rect -1580 317 -1498 355
rect -1580 283 -1556 317
rect -1522 283 -1498 317
rect -1580 245 -1498 283
rect -1580 211 -1556 245
rect -1522 211 -1498 245
rect -1580 173 -1498 211
rect -1580 139 -1556 173
rect -1522 139 -1498 173
rect -1580 101 -1498 139
rect -1580 67 -1556 101
rect -1522 67 -1498 101
rect -1580 29 -1498 67
rect -1580 -5 -1556 29
rect -1522 -5 -1498 29
rect -1580 -43 -1498 -5
rect -1580 -77 -1556 -43
rect -1522 -77 -1498 -43
rect -1580 -115 -1498 -77
rect -1580 -149 -1556 -115
rect -1522 -149 -1498 -115
rect -1580 -187 -1498 -149
rect -1580 -221 -1556 -187
rect -1522 -221 -1498 -187
rect -1580 -259 -1498 -221
rect -1580 -293 -1556 -259
rect -1522 -293 -1498 -259
rect -1580 -331 -1498 -293
rect -1580 -365 -1556 -331
rect -1522 -365 -1498 -331
rect -1580 -403 -1498 -365
rect -1580 -437 -1556 -403
rect -1522 -437 -1498 -403
rect -1580 -475 -1498 -437
rect -1580 -509 -1556 -475
rect -1522 -509 -1498 -475
rect -1580 -547 -1498 -509
rect -1580 -581 -1556 -547
rect -1522 -581 -1498 -547
rect -1580 -619 -1498 -581
rect -1580 -653 -1556 -619
rect -1522 -653 -1498 -619
rect -1580 -691 -1498 -653
rect -1580 -725 -1556 -691
rect -1522 -725 -1498 -691
rect -1580 -763 -1498 -725
rect -1580 -797 -1556 -763
rect -1522 -797 -1498 -763
rect -1580 -835 -1498 -797
rect -1580 -869 -1556 -835
rect -1522 -869 -1498 -835
rect -1580 -907 -1498 -869
rect -1580 -941 -1556 -907
rect -1522 -941 -1498 -907
rect -1580 -979 -1498 -941
rect -1580 -1013 -1556 -979
rect -1522 -1013 -1498 -979
rect -1580 -1051 -1498 -1013
rect -798 6998 948 7022
rect -798 6820 -554 6998
rect 704 6820 948 6998
rect -798 6757 948 6820
rect -798 6650 -716 6757
rect -798 6616 -774 6650
rect -740 6616 -716 6650
rect -798 6578 -716 6616
rect -798 6544 -774 6578
rect -740 6544 -716 6578
rect -798 6506 -716 6544
rect -798 6472 -774 6506
rect -740 6472 -716 6506
rect -798 6434 -716 6472
rect -798 6400 -774 6434
rect -740 6400 -716 6434
rect -798 6362 -716 6400
rect -798 6328 -774 6362
rect -740 6328 -716 6362
rect -798 6290 -716 6328
rect -798 6256 -774 6290
rect -740 6256 -716 6290
rect -798 6218 -716 6256
rect -798 6184 -774 6218
rect -740 6184 -716 6218
rect -798 6146 -716 6184
rect 866 6650 948 6757
rect 866 6616 890 6650
rect 924 6616 948 6650
rect 866 6578 948 6616
rect 866 6544 890 6578
rect 924 6544 948 6578
rect 866 6506 948 6544
rect 866 6472 890 6506
rect 924 6472 948 6506
rect 866 6434 948 6472
rect 866 6400 890 6434
rect 924 6400 948 6434
rect 866 6362 948 6400
rect 866 6328 890 6362
rect 924 6328 948 6362
rect 866 6290 948 6328
rect 866 6256 890 6290
rect 924 6256 948 6290
rect 866 6218 948 6256
rect 866 6184 890 6218
rect 924 6184 948 6218
rect -798 6112 -774 6146
rect -740 6112 -716 6146
rect -798 6074 -716 6112
rect -798 6040 -774 6074
rect -740 6040 -716 6074
rect -798 6002 -716 6040
rect -798 5968 -774 6002
rect -740 5968 -716 6002
rect -798 5930 -716 5968
rect -798 5896 -774 5930
rect -740 5896 -716 5930
rect -798 5858 -716 5896
rect -798 5824 -774 5858
rect -740 5824 -716 5858
rect -798 5786 -716 5824
rect -798 5752 -774 5786
rect -740 5752 -716 5786
rect -798 5714 -716 5752
rect -798 5680 -774 5714
rect -740 5680 -716 5714
rect -798 5642 -716 5680
rect -798 5608 -774 5642
rect -740 5608 -716 5642
rect -798 5570 -716 5608
rect -798 5536 -774 5570
rect -740 5536 -716 5570
rect -798 5498 -716 5536
rect -798 5464 -774 5498
rect -740 5464 -716 5498
rect -798 5426 -716 5464
rect -798 5392 -774 5426
rect -740 5392 -716 5426
rect -798 5354 -716 5392
rect -798 5320 -774 5354
rect -740 5320 -716 5354
rect -798 5282 -716 5320
rect -798 5248 -774 5282
rect -740 5248 -716 5282
rect -798 5210 -716 5248
rect -798 5176 -774 5210
rect -740 5176 -716 5210
rect -798 5138 -716 5176
rect -798 5104 -774 5138
rect -740 5104 -716 5138
rect -798 5066 -716 5104
rect -798 5032 -774 5066
rect -740 5032 -716 5066
rect -798 4994 -716 5032
rect -798 4960 -774 4994
rect -740 4960 -716 4994
rect -798 4922 -716 4960
rect -798 4888 -774 4922
rect -740 4888 -716 4922
rect -798 4850 -716 4888
rect -798 4816 -774 4850
rect -740 4816 -716 4850
rect -798 4778 -716 4816
rect -798 4744 -774 4778
rect -740 4744 -716 4778
rect -798 4706 -716 4744
rect -798 4672 -774 4706
rect -740 4672 -716 4706
rect -798 4634 -716 4672
rect -798 4600 -774 4634
rect -740 4600 -716 4634
rect -798 4562 -716 4600
rect -798 4528 -774 4562
rect -740 4528 -716 4562
rect -798 4490 -716 4528
rect -798 4456 -774 4490
rect -740 4456 -716 4490
rect -798 4418 -716 4456
rect -798 4384 -774 4418
rect -740 4384 -716 4418
rect -798 4346 -716 4384
rect -798 4312 -774 4346
rect -740 4312 -716 4346
rect -798 4274 -716 4312
rect -798 4240 -774 4274
rect -740 4240 -716 4274
rect -798 4202 -716 4240
rect -798 4168 -774 4202
rect -740 4168 -716 4202
rect -798 4130 -716 4168
rect -798 4096 -774 4130
rect -740 4096 -716 4130
rect -798 4058 -716 4096
rect -798 4024 -774 4058
rect -740 4024 -716 4058
rect -798 3986 -716 4024
rect -798 3952 -774 3986
rect -740 3952 -716 3986
rect -798 3914 -716 3952
rect -798 3880 -774 3914
rect -740 3880 -716 3914
rect -798 3842 -716 3880
rect -798 3808 -774 3842
rect -740 3808 -716 3842
rect -798 3770 -716 3808
rect -798 3736 -774 3770
rect -740 3736 -716 3770
rect -798 3698 -716 3736
rect -798 3664 -774 3698
rect -740 3664 -716 3698
rect -798 3626 -716 3664
rect -798 3592 -774 3626
rect -740 3592 -716 3626
rect -798 3554 -716 3592
rect -798 3520 -774 3554
rect -740 3520 -716 3554
rect -798 3482 -716 3520
rect -798 3448 -774 3482
rect -740 3448 -716 3482
rect -798 3410 -716 3448
rect -798 3376 -774 3410
rect -740 3376 -716 3410
rect -798 3338 -716 3376
rect -798 3304 -774 3338
rect -740 3304 -716 3338
rect -798 3266 -716 3304
rect -798 3232 -774 3266
rect -740 3232 -716 3266
rect -798 3194 -716 3232
rect -798 3160 -774 3194
rect -740 3160 -716 3194
rect -798 3122 -716 3160
rect -798 3088 -774 3122
rect -740 3088 -716 3122
rect -798 3050 -716 3088
rect -798 3016 -774 3050
rect -740 3016 -716 3050
rect -798 2978 -716 3016
rect -798 2944 -774 2978
rect -740 2944 -716 2978
rect -798 2906 -716 2944
rect -798 2872 -774 2906
rect -740 2872 -716 2906
rect -798 2834 -716 2872
rect -798 2800 -774 2834
rect -740 2800 -716 2834
rect -798 2762 -716 2800
rect -798 2728 -774 2762
rect -740 2728 -716 2762
rect -798 2690 -716 2728
rect -798 2656 -774 2690
rect -740 2656 -716 2690
rect -798 2618 -716 2656
rect -798 2584 -774 2618
rect -740 2584 -716 2618
rect -798 2546 -716 2584
rect -798 2512 -774 2546
rect -740 2512 -716 2546
rect -798 2474 -716 2512
rect -798 2440 -774 2474
rect -740 2440 -716 2474
rect -798 2402 -716 2440
rect -798 2368 -774 2402
rect -740 2368 -716 2402
rect -798 2330 -716 2368
rect -798 2296 -774 2330
rect -740 2296 -716 2330
rect -798 2258 -716 2296
rect -798 2224 -774 2258
rect -740 2224 -716 2258
rect -798 2186 -716 2224
rect -798 2152 -774 2186
rect -740 2152 -716 2186
rect -798 2114 -716 2152
rect -798 2080 -774 2114
rect -740 2080 -716 2114
rect -798 2042 -716 2080
rect -798 2008 -774 2042
rect -740 2008 -716 2042
rect -798 1970 -716 2008
rect -798 1936 -774 1970
rect -740 1936 -716 1970
rect -798 1898 -716 1936
rect -798 1864 -774 1898
rect -740 1864 -716 1898
rect -798 1826 -716 1864
rect -798 1792 -774 1826
rect -740 1792 -716 1826
rect -798 1754 -716 1792
rect -798 1720 -774 1754
rect -740 1720 -716 1754
rect -798 1682 -716 1720
rect -798 1648 -774 1682
rect -740 1648 -716 1682
rect -798 1610 -716 1648
rect -798 1576 -774 1610
rect -740 1576 -716 1610
rect -798 1538 -716 1576
rect -798 1504 -774 1538
rect -740 1504 -716 1538
rect -798 1466 -716 1504
rect -798 1432 -774 1466
rect -740 1432 -716 1466
rect -798 1394 -716 1432
rect -798 1360 -774 1394
rect -740 1360 -716 1394
rect -798 1322 -716 1360
rect -798 1288 -774 1322
rect -740 1288 -716 1322
rect -798 1250 -716 1288
rect -798 1216 -774 1250
rect -740 1216 -716 1250
rect -798 1178 -716 1216
rect -798 1144 -774 1178
rect -740 1144 -716 1178
rect -798 1106 -716 1144
rect -798 1072 -774 1106
rect -740 1072 -716 1106
rect -798 1034 -716 1072
rect -798 1000 -774 1034
rect -740 1000 -716 1034
rect -798 962 -716 1000
rect -798 928 -774 962
rect -740 928 -716 962
rect -798 890 -716 928
rect -798 856 -774 890
rect -740 856 -716 890
rect -798 818 -716 856
rect -798 784 -774 818
rect -740 784 -716 818
rect -798 746 -716 784
rect -798 712 -774 746
rect -740 712 -716 746
rect -798 674 -716 712
rect -798 640 -774 674
rect -740 640 -716 674
rect -798 602 -716 640
rect -798 568 -774 602
rect -740 568 -716 602
rect -798 530 -716 568
rect -798 496 -774 530
rect -740 496 -716 530
rect -798 458 -716 496
rect -798 424 -774 458
rect -740 424 -716 458
rect -798 386 -716 424
rect -798 352 -774 386
rect -740 352 -716 386
rect -798 314 -716 352
rect -798 280 -774 314
rect -740 280 -716 314
rect -798 242 -716 280
rect -798 208 -774 242
rect -740 208 -716 242
rect -798 170 -716 208
rect -798 136 -774 170
rect -740 136 -716 170
rect -798 98 -716 136
rect -798 64 -774 98
rect -740 64 -716 98
rect -798 26 -716 64
rect -798 -8 -774 26
rect -740 -8 -716 26
rect -798 -46 -716 -8
rect -798 -80 -774 -46
rect -740 -80 -716 -46
rect -798 -118 -716 -80
rect -798 -152 -774 -118
rect -740 -152 -716 -118
rect -798 -190 -716 -152
rect -659 6146 -457 6165
rect -659 -152 -647 6146
rect -469 -152 -457 6146
rect -659 -164 -457 -152
rect -134 6146 284 6165
rect -134 -152 -122 6146
rect 272 -152 284 6146
rect -134 -164 284 -152
rect 607 6146 809 6165
rect 607 -152 619 6146
rect 797 -152 809 6146
rect 607 -164 809 -152
rect 866 6146 948 6184
rect 866 6112 890 6146
rect 924 6112 948 6146
rect 866 6074 948 6112
rect 866 6040 890 6074
rect 924 6040 948 6074
rect 866 6002 948 6040
rect 866 5968 890 6002
rect 924 5968 948 6002
rect 866 5930 948 5968
rect 866 5896 890 5930
rect 924 5896 948 5930
rect 866 5858 948 5896
rect 866 5824 890 5858
rect 924 5824 948 5858
rect 866 5786 948 5824
rect 866 5752 890 5786
rect 924 5752 948 5786
rect 866 5714 948 5752
rect 866 5680 890 5714
rect 924 5680 948 5714
rect 866 5642 948 5680
rect 866 5608 890 5642
rect 924 5608 948 5642
rect 866 5570 948 5608
rect 866 5536 890 5570
rect 924 5536 948 5570
rect 866 5498 948 5536
rect 866 5464 890 5498
rect 924 5464 948 5498
rect 866 5426 948 5464
rect 866 5392 890 5426
rect 924 5392 948 5426
rect 866 5354 948 5392
rect 866 5320 890 5354
rect 924 5320 948 5354
rect 866 5282 948 5320
rect 866 5248 890 5282
rect 924 5248 948 5282
rect 866 5210 948 5248
rect 866 5176 890 5210
rect 924 5176 948 5210
rect 866 5138 948 5176
rect 866 5104 890 5138
rect 924 5104 948 5138
rect 866 5066 948 5104
rect 866 5032 890 5066
rect 924 5032 948 5066
rect 866 4994 948 5032
rect 866 4960 890 4994
rect 924 4960 948 4994
rect 866 4922 948 4960
rect 866 4888 890 4922
rect 924 4888 948 4922
rect 866 4850 948 4888
rect 866 4816 890 4850
rect 924 4816 948 4850
rect 866 4778 948 4816
rect 866 4744 890 4778
rect 924 4744 948 4778
rect 866 4706 948 4744
rect 866 4672 890 4706
rect 924 4672 948 4706
rect 866 4634 948 4672
rect 866 4600 890 4634
rect 924 4600 948 4634
rect 866 4562 948 4600
rect 866 4528 890 4562
rect 924 4528 948 4562
rect 866 4490 948 4528
rect 866 4456 890 4490
rect 924 4456 948 4490
rect 866 4418 948 4456
rect 866 4384 890 4418
rect 924 4384 948 4418
rect 866 4346 948 4384
rect 866 4312 890 4346
rect 924 4312 948 4346
rect 866 4274 948 4312
rect 866 4240 890 4274
rect 924 4240 948 4274
rect 866 4202 948 4240
rect 866 4168 890 4202
rect 924 4168 948 4202
rect 866 4130 948 4168
rect 866 4096 890 4130
rect 924 4096 948 4130
rect 866 4058 948 4096
rect 866 4024 890 4058
rect 924 4024 948 4058
rect 866 3986 948 4024
rect 866 3952 890 3986
rect 924 3952 948 3986
rect 866 3914 948 3952
rect 866 3880 890 3914
rect 924 3880 948 3914
rect 866 3842 948 3880
rect 866 3808 890 3842
rect 924 3808 948 3842
rect 866 3770 948 3808
rect 866 3736 890 3770
rect 924 3736 948 3770
rect 866 3698 948 3736
rect 866 3664 890 3698
rect 924 3664 948 3698
rect 866 3626 948 3664
rect 866 3592 890 3626
rect 924 3592 948 3626
rect 866 3554 948 3592
rect 866 3520 890 3554
rect 924 3520 948 3554
rect 866 3482 948 3520
rect 866 3448 890 3482
rect 924 3448 948 3482
rect 866 3410 948 3448
rect 866 3376 890 3410
rect 924 3376 948 3410
rect 866 3338 948 3376
rect 866 3304 890 3338
rect 924 3304 948 3338
rect 866 3266 948 3304
rect 866 3232 890 3266
rect 924 3232 948 3266
rect 866 3194 948 3232
rect 866 3160 890 3194
rect 924 3160 948 3194
rect 866 3122 948 3160
rect 866 3088 890 3122
rect 924 3088 948 3122
rect 866 3050 948 3088
rect 866 3016 890 3050
rect 924 3016 948 3050
rect 866 2978 948 3016
rect 866 2944 890 2978
rect 924 2944 948 2978
rect 866 2906 948 2944
rect 866 2872 890 2906
rect 924 2872 948 2906
rect 866 2834 948 2872
rect 866 2800 890 2834
rect 924 2800 948 2834
rect 866 2762 948 2800
rect 866 2728 890 2762
rect 924 2728 948 2762
rect 866 2690 948 2728
rect 866 2656 890 2690
rect 924 2656 948 2690
rect 866 2618 948 2656
rect 866 2584 890 2618
rect 924 2584 948 2618
rect 866 2546 948 2584
rect 866 2512 890 2546
rect 924 2512 948 2546
rect 866 2474 948 2512
rect 866 2440 890 2474
rect 924 2440 948 2474
rect 866 2402 948 2440
rect 866 2368 890 2402
rect 924 2368 948 2402
rect 866 2330 948 2368
rect 866 2296 890 2330
rect 924 2296 948 2330
rect 866 2258 948 2296
rect 866 2224 890 2258
rect 924 2224 948 2258
rect 866 2186 948 2224
rect 866 2152 890 2186
rect 924 2152 948 2186
rect 866 2114 948 2152
rect 866 2080 890 2114
rect 924 2080 948 2114
rect 866 2042 948 2080
rect 866 2008 890 2042
rect 924 2008 948 2042
rect 866 1970 948 2008
rect 866 1936 890 1970
rect 924 1936 948 1970
rect 866 1898 948 1936
rect 866 1864 890 1898
rect 924 1864 948 1898
rect 866 1826 948 1864
rect 866 1792 890 1826
rect 924 1792 948 1826
rect 866 1754 948 1792
rect 866 1720 890 1754
rect 924 1720 948 1754
rect 866 1682 948 1720
rect 866 1648 890 1682
rect 924 1648 948 1682
rect 866 1610 948 1648
rect 866 1576 890 1610
rect 924 1576 948 1610
rect 866 1538 948 1576
rect 866 1504 890 1538
rect 924 1504 948 1538
rect 866 1466 948 1504
rect 866 1432 890 1466
rect 924 1432 948 1466
rect 866 1394 948 1432
rect 866 1360 890 1394
rect 924 1360 948 1394
rect 866 1322 948 1360
rect 866 1288 890 1322
rect 924 1288 948 1322
rect 866 1250 948 1288
rect 866 1216 890 1250
rect 924 1216 948 1250
rect 866 1178 948 1216
rect 866 1144 890 1178
rect 924 1144 948 1178
rect 866 1106 948 1144
rect 866 1072 890 1106
rect 924 1072 948 1106
rect 866 1034 948 1072
rect 866 1000 890 1034
rect 924 1000 948 1034
rect 866 962 948 1000
rect 866 928 890 962
rect 924 928 948 962
rect 866 890 948 928
rect 866 856 890 890
rect 924 856 948 890
rect 866 818 948 856
rect 866 784 890 818
rect 924 784 948 818
rect 866 746 948 784
rect 866 712 890 746
rect 924 712 948 746
rect 866 674 948 712
rect 866 640 890 674
rect 924 640 948 674
rect 866 602 948 640
rect 866 568 890 602
rect 924 568 948 602
rect 866 530 948 568
rect 866 496 890 530
rect 924 496 948 530
rect 866 458 948 496
rect 866 424 890 458
rect 924 424 948 458
rect 866 386 948 424
rect 866 352 890 386
rect 924 352 948 386
rect 866 314 948 352
rect 866 280 890 314
rect 924 280 948 314
rect 866 242 948 280
rect 866 208 890 242
rect 924 208 948 242
rect 866 170 948 208
rect 866 136 890 170
rect 924 136 948 170
rect 866 98 948 136
rect 866 64 890 98
rect 924 64 948 98
rect 866 26 948 64
rect 866 -8 890 26
rect 924 -8 948 26
rect 866 -46 948 -8
rect 866 -80 890 -46
rect 924 -80 948 -46
rect 866 -118 948 -80
rect 866 -152 890 -118
rect 924 -152 948 -118
rect -798 -224 -774 -190
rect -740 -224 -716 -190
rect -798 -262 -716 -224
rect -798 -296 -774 -262
rect -740 -296 -716 -262
rect -798 -334 -716 -296
rect -798 -368 -774 -334
rect -740 -368 -716 -334
rect -798 -406 -716 -368
rect -798 -440 -774 -406
rect -740 -440 -716 -406
rect -798 -478 -716 -440
rect 866 -190 948 -152
rect 866 -224 890 -190
rect 924 -224 948 -190
rect 866 -262 948 -224
rect 866 -296 890 -262
rect 924 -296 948 -262
rect 866 -334 948 -296
rect 866 -368 890 -334
rect 924 -368 948 -334
rect 866 -406 948 -368
rect 866 -440 890 -406
rect 924 -440 948 -406
rect -798 -512 -774 -478
rect -740 -512 -716 -478
rect -798 -550 -716 -512
rect -798 -584 -774 -550
rect -740 -584 -716 -550
rect -798 -622 -716 -584
rect -798 -656 -774 -622
rect -740 -656 -716 -622
rect -798 -757 -716 -656
rect -146 -459 290 -443
rect -146 -493 -130 -459
rect -96 -493 -56 -459
rect -22 -493 18 -459
rect 52 -493 92 -459
rect 126 -493 166 -459
rect 200 -493 240 -459
rect 274 -493 290 -459
rect -146 -533 290 -493
rect -146 -567 -130 -533
rect -96 -567 -56 -533
rect -22 -567 18 -533
rect 52 -567 92 -533
rect 126 -567 166 -533
rect 200 -567 240 -533
rect 274 -567 290 -533
rect -146 -607 290 -567
rect -146 -641 -130 -607
rect -96 -641 -56 -607
rect -22 -641 18 -607
rect 52 -641 92 -607
rect 126 -641 166 -607
rect 200 -641 240 -607
rect 274 -641 290 -607
rect -146 -657 290 -641
rect 866 -478 948 -440
rect 866 -512 890 -478
rect 924 -512 948 -478
rect 866 -550 948 -512
rect 866 -584 890 -550
rect 924 -584 948 -550
rect 866 -622 948 -584
rect 866 -656 890 -622
rect 924 -656 948 -622
rect 866 -757 948 -656
rect -798 -820 948 -757
rect -798 -998 -554 -820
rect 704 -998 948 -820
rect -798 -1022 948 -998
rect 1648 7013 1730 7051
rect 1648 6979 1672 7013
rect 1706 6979 1730 7013
rect 1648 6941 1730 6979
rect 1648 6907 1672 6941
rect 1706 6907 1730 6941
rect 1648 6869 1730 6907
rect 1648 6835 1672 6869
rect 1706 6835 1730 6869
rect 1648 6797 1730 6835
rect 1648 6763 1672 6797
rect 1706 6763 1730 6797
rect 1648 6725 1730 6763
rect 1648 6691 1672 6725
rect 1706 6691 1730 6725
rect 1648 6653 1730 6691
rect 1648 6619 1672 6653
rect 1706 6619 1730 6653
rect 1648 6581 1730 6619
rect 1648 6547 1672 6581
rect 1706 6547 1730 6581
rect 1648 6509 1730 6547
rect 1648 6475 1672 6509
rect 1706 6475 1730 6509
rect 1648 6437 1730 6475
rect 1648 6403 1672 6437
rect 1706 6403 1730 6437
rect 1648 6365 1730 6403
rect 1648 6331 1672 6365
rect 1706 6331 1730 6365
rect 1648 6293 1730 6331
rect 1648 6259 1672 6293
rect 1706 6259 1730 6293
rect 1648 6221 1730 6259
rect 1648 6187 1672 6221
rect 1706 6187 1730 6221
rect 1648 6149 1730 6187
rect 1648 6115 1672 6149
rect 1706 6115 1730 6149
rect 1648 6077 1730 6115
rect 1648 6043 1672 6077
rect 1706 6043 1730 6077
rect 1648 6005 1730 6043
rect 1648 5971 1672 6005
rect 1706 5971 1730 6005
rect 1648 5933 1730 5971
rect 1648 5899 1672 5933
rect 1706 5899 1730 5933
rect 1648 5861 1730 5899
rect 1648 5827 1672 5861
rect 1706 5827 1730 5861
rect 1648 5789 1730 5827
rect 1648 5755 1672 5789
rect 1706 5755 1730 5789
rect 1648 5717 1730 5755
rect 1648 5683 1672 5717
rect 1706 5683 1730 5717
rect 1648 5645 1730 5683
rect 1648 5611 1672 5645
rect 1706 5611 1730 5645
rect 1648 5573 1730 5611
rect 1648 5539 1672 5573
rect 1706 5539 1730 5573
rect 1648 5501 1730 5539
rect 1648 5467 1672 5501
rect 1706 5467 1730 5501
rect 1648 5429 1730 5467
rect 1648 5395 1672 5429
rect 1706 5395 1730 5429
rect 1648 5357 1730 5395
rect 1648 5323 1672 5357
rect 1706 5323 1730 5357
rect 1648 5285 1730 5323
rect 1648 5251 1672 5285
rect 1706 5251 1730 5285
rect 1648 5213 1730 5251
rect 1648 5179 1672 5213
rect 1706 5179 1730 5213
rect 1648 5141 1730 5179
rect 1648 5107 1672 5141
rect 1706 5107 1730 5141
rect 1648 5069 1730 5107
rect 1648 5035 1672 5069
rect 1706 5035 1730 5069
rect 1648 4997 1730 5035
rect 1648 4963 1672 4997
rect 1706 4963 1730 4997
rect 1648 4925 1730 4963
rect 1648 4891 1672 4925
rect 1706 4891 1730 4925
rect 1648 4853 1730 4891
rect 1648 4819 1672 4853
rect 1706 4819 1730 4853
rect 1648 4781 1730 4819
rect 1648 4747 1672 4781
rect 1706 4747 1730 4781
rect 1648 4709 1730 4747
rect 1648 4675 1672 4709
rect 1706 4675 1730 4709
rect 1648 4637 1730 4675
rect 1648 4603 1672 4637
rect 1706 4603 1730 4637
rect 1648 4565 1730 4603
rect 1648 4531 1672 4565
rect 1706 4531 1730 4565
rect 1648 4493 1730 4531
rect 1648 4459 1672 4493
rect 1706 4459 1730 4493
rect 1648 4421 1730 4459
rect 1648 4387 1672 4421
rect 1706 4387 1730 4421
rect 1648 4349 1730 4387
rect 1648 4315 1672 4349
rect 1706 4315 1730 4349
rect 1648 4277 1730 4315
rect 1648 4243 1672 4277
rect 1706 4243 1730 4277
rect 1648 4205 1730 4243
rect 1648 4171 1672 4205
rect 1706 4171 1730 4205
rect 1648 4133 1730 4171
rect 1648 4099 1672 4133
rect 1706 4099 1730 4133
rect 1648 4061 1730 4099
rect 1648 4027 1672 4061
rect 1706 4027 1730 4061
rect 1648 3989 1730 4027
rect 1648 3955 1672 3989
rect 1706 3955 1730 3989
rect 1648 3917 1730 3955
rect 1648 3883 1672 3917
rect 1706 3883 1730 3917
rect 1648 3845 1730 3883
rect 1648 3811 1672 3845
rect 1706 3811 1730 3845
rect 1648 3773 1730 3811
rect 1648 3739 1672 3773
rect 1706 3739 1730 3773
rect 1648 3701 1730 3739
rect 1648 3667 1672 3701
rect 1706 3667 1730 3701
rect 1648 3629 1730 3667
rect 1648 3595 1672 3629
rect 1706 3595 1730 3629
rect 1648 3557 1730 3595
rect 1648 3523 1672 3557
rect 1706 3523 1730 3557
rect 1648 3485 1730 3523
rect 1648 3451 1672 3485
rect 1706 3451 1730 3485
rect 1648 3413 1730 3451
rect 1648 3379 1672 3413
rect 1706 3379 1730 3413
rect 1648 3341 1730 3379
rect 1648 3307 1672 3341
rect 1706 3307 1730 3341
rect 1648 3269 1730 3307
rect 1648 3235 1672 3269
rect 1706 3235 1730 3269
rect 1648 3197 1730 3235
rect 1648 3163 1672 3197
rect 1706 3163 1730 3197
rect 1648 3125 1730 3163
rect 1648 3091 1672 3125
rect 1706 3091 1730 3125
rect 1648 3053 1730 3091
rect 1648 3019 1672 3053
rect 1706 3019 1730 3053
rect 1648 2981 1730 3019
rect 1648 2947 1672 2981
rect 1706 2947 1730 2981
rect 1648 2909 1730 2947
rect 1648 2875 1672 2909
rect 1706 2875 1730 2909
rect 1648 2837 1730 2875
rect 1648 2803 1672 2837
rect 1706 2803 1730 2837
rect 1648 2765 1730 2803
rect 1648 2731 1672 2765
rect 1706 2731 1730 2765
rect 1648 2693 1730 2731
rect 1648 2659 1672 2693
rect 1706 2659 1730 2693
rect 1648 2621 1730 2659
rect 1648 2587 1672 2621
rect 1706 2587 1730 2621
rect 1648 2549 1730 2587
rect 1648 2515 1672 2549
rect 1706 2515 1730 2549
rect 1648 2477 1730 2515
rect 1648 2443 1672 2477
rect 1706 2443 1730 2477
rect 1648 2405 1730 2443
rect 1648 2371 1672 2405
rect 1706 2371 1730 2405
rect 1648 2333 1730 2371
rect 1648 2299 1672 2333
rect 1706 2299 1730 2333
rect 1648 2261 1730 2299
rect 1648 2227 1672 2261
rect 1706 2227 1730 2261
rect 1648 2189 1730 2227
rect 1648 2155 1672 2189
rect 1706 2155 1730 2189
rect 1648 2117 1730 2155
rect 1648 2083 1672 2117
rect 1706 2083 1730 2117
rect 1648 2045 1730 2083
rect 1648 2011 1672 2045
rect 1706 2011 1730 2045
rect 1648 1973 1730 2011
rect 1648 1939 1672 1973
rect 1706 1939 1730 1973
rect 1648 1901 1730 1939
rect 1648 1867 1672 1901
rect 1706 1867 1730 1901
rect 1648 1829 1730 1867
rect 1648 1795 1672 1829
rect 1706 1795 1730 1829
rect 1648 1757 1730 1795
rect 1648 1723 1672 1757
rect 1706 1723 1730 1757
rect 1648 1685 1730 1723
rect 1648 1651 1672 1685
rect 1706 1651 1730 1685
rect 1648 1613 1730 1651
rect 1648 1579 1672 1613
rect 1706 1579 1730 1613
rect 1648 1541 1730 1579
rect 1648 1507 1672 1541
rect 1706 1507 1730 1541
rect 1648 1469 1730 1507
rect 1648 1435 1672 1469
rect 1706 1435 1730 1469
rect 1648 1397 1730 1435
rect 1648 1363 1672 1397
rect 1706 1363 1730 1397
rect 1648 1325 1730 1363
rect 1648 1291 1672 1325
rect 1706 1291 1730 1325
rect 1648 1253 1730 1291
rect 1648 1219 1672 1253
rect 1706 1219 1730 1253
rect 1648 1181 1730 1219
rect 1648 1147 1672 1181
rect 1706 1147 1730 1181
rect 1648 1109 1730 1147
rect 1648 1075 1672 1109
rect 1706 1075 1730 1109
rect 1648 1037 1730 1075
rect 1648 1003 1672 1037
rect 1706 1003 1730 1037
rect 1648 965 1730 1003
rect 1648 931 1672 965
rect 1706 931 1730 965
rect 1648 893 1730 931
rect 1648 859 1672 893
rect 1706 859 1730 893
rect 1648 821 1730 859
rect 1648 787 1672 821
rect 1706 787 1730 821
rect 1648 749 1730 787
rect 1648 715 1672 749
rect 1706 715 1730 749
rect 1648 677 1730 715
rect 1648 643 1672 677
rect 1706 643 1730 677
rect 1648 605 1730 643
rect 1648 571 1672 605
rect 1706 571 1730 605
rect 1648 533 1730 571
rect 1648 499 1672 533
rect 1706 499 1730 533
rect 1648 461 1730 499
rect 1648 427 1672 461
rect 1706 427 1730 461
rect 1648 389 1730 427
rect 1648 355 1672 389
rect 1706 355 1730 389
rect 1648 317 1730 355
rect 1648 283 1672 317
rect 1706 283 1730 317
rect 1648 245 1730 283
rect 1648 211 1672 245
rect 1706 211 1730 245
rect 1648 173 1730 211
rect 1648 139 1672 173
rect 1706 139 1730 173
rect 1648 101 1730 139
rect 1648 67 1672 101
rect 1706 67 1730 101
rect 1648 29 1730 67
rect 1648 -5 1672 29
rect 1706 -5 1730 29
rect 1648 -43 1730 -5
rect 1648 -77 1672 -43
rect 1706 -77 1730 -43
rect 1648 -115 1730 -77
rect 1648 -149 1672 -115
rect 1706 -149 1730 -115
rect 1648 -187 1730 -149
rect 1648 -221 1672 -187
rect 1706 -221 1730 -187
rect 1648 -259 1730 -221
rect 1648 -293 1672 -259
rect 1706 -293 1730 -259
rect 1648 -331 1730 -293
rect 1648 -365 1672 -331
rect 1706 -365 1730 -331
rect 1648 -403 1730 -365
rect 1648 -437 1672 -403
rect 1706 -437 1730 -403
rect 1648 -475 1730 -437
rect 1648 -509 1672 -475
rect 1706 -509 1730 -475
rect 1648 -547 1730 -509
rect 1648 -581 1672 -547
rect 1706 -581 1730 -547
rect 1648 -619 1730 -581
rect 1648 -653 1672 -619
rect 1706 -653 1730 -619
rect 1648 -691 1730 -653
rect 1648 -725 1672 -691
rect 1706 -725 1730 -691
rect 1648 -763 1730 -725
rect 1648 -797 1672 -763
rect 1706 -797 1730 -763
rect 1648 -835 1730 -797
rect 1648 -869 1672 -835
rect 1706 -869 1730 -835
rect 1648 -907 1730 -869
rect 1648 -941 1672 -907
rect 1706 -941 1730 -907
rect 1648 -979 1730 -941
rect 1648 -1013 1672 -979
rect 1706 -1013 1730 -979
rect -1580 -1085 -1556 -1051
rect -1522 -1085 -1498 -1051
rect -1580 -1123 -1498 -1085
rect -1580 -1157 -1556 -1123
rect -1522 -1157 -1498 -1123
rect -1580 -1195 -1498 -1157
rect -1580 -1229 -1556 -1195
rect -1522 -1229 -1498 -1195
rect -1580 -1267 -1498 -1229
rect -1580 -1301 -1556 -1267
rect -1522 -1301 -1498 -1267
rect -1580 -1339 -1498 -1301
rect -1580 -1373 -1556 -1339
rect -1522 -1373 -1498 -1339
rect -1580 -1411 -1498 -1373
rect -1580 -1445 -1556 -1411
rect -1522 -1445 -1498 -1411
rect -1580 -1483 -1498 -1445
rect -1580 -1517 -1556 -1483
rect -1522 -1517 -1498 -1483
rect -1580 -1555 -1498 -1517
rect -1580 -1589 -1556 -1555
rect -1522 -1589 -1498 -1555
rect -1580 -1627 -1498 -1589
rect -1580 -1661 -1556 -1627
rect -1522 -1661 -1498 -1627
rect -1580 -1722 -1498 -1661
rect 1648 -1051 1730 -1013
rect 1648 -1085 1672 -1051
rect 1706 -1085 1730 -1051
rect 1648 -1123 1730 -1085
rect 1648 -1157 1672 -1123
rect 1706 -1157 1730 -1123
rect 1648 -1195 1730 -1157
rect 1648 -1229 1672 -1195
rect 1706 -1229 1730 -1195
rect 1648 -1267 1730 -1229
rect 1648 -1301 1672 -1267
rect 1706 -1301 1730 -1267
rect 1648 -1339 1730 -1301
rect 1648 -1373 1672 -1339
rect 1706 -1373 1730 -1339
rect 1648 -1411 1730 -1373
rect 1648 -1445 1672 -1411
rect 1706 -1445 1730 -1411
rect 1648 -1483 1730 -1445
rect 1648 -1517 1672 -1483
rect 1706 -1517 1730 -1483
rect 1648 -1555 1730 -1517
rect 1648 -1589 1672 -1555
rect 1706 -1589 1730 -1555
rect 1648 -1627 1730 -1589
rect 1648 -1661 1672 -1627
rect 1706 -1661 1730 -1627
rect 1648 -1722 1730 -1661
rect -1580 -1746 1730 -1722
rect -1580 -1780 -1454 -1746
rect -1420 -1780 -1382 -1746
rect -1348 -1780 -1310 -1746
rect -1276 -1780 -1238 -1746
rect -1204 -1780 -1166 -1746
rect -1132 -1780 -1094 -1746
rect -1060 -1780 -1022 -1746
rect -988 -1780 -950 -1746
rect -916 -1780 -878 -1746
rect -844 -1780 -806 -1746
rect -772 -1780 -734 -1746
rect -700 -1780 -662 -1746
rect -628 -1780 -590 -1746
rect -556 -1780 -518 -1746
rect -484 -1780 -446 -1746
rect -412 -1780 -374 -1746
rect -340 -1780 -302 -1746
rect -268 -1780 -230 -1746
rect -196 -1780 -158 -1746
rect -124 -1780 -86 -1746
rect -52 -1780 -14 -1746
rect 20 -1780 58 -1746
rect 92 -1780 130 -1746
rect 164 -1780 202 -1746
rect 236 -1780 274 -1746
rect 308 -1780 346 -1746
rect 380 -1780 418 -1746
rect 452 -1780 490 -1746
rect 524 -1780 562 -1746
rect 596 -1780 634 -1746
rect 668 -1780 706 -1746
rect 740 -1780 778 -1746
rect 812 -1780 850 -1746
rect 884 -1780 922 -1746
rect 956 -1780 994 -1746
rect 1028 -1780 1066 -1746
rect 1100 -1780 1138 -1746
rect 1172 -1780 1210 -1746
rect 1244 -1780 1282 -1746
rect 1316 -1780 1354 -1746
rect 1388 -1780 1426 -1746
rect 1460 -1780 1498 -1746
rect 1532 -1780 1570 -1746
rect 1604 -1780 1730 -1746
rect -1580 -1804 1730 -1780
<< viali >>
rect -1454 7746 -1420 7780
rect -1382 7746 -1348 7780
rect -1310 7746 -1276 7780
rect -1238 7746 -1204 7780
rect -1166 7746 -1132 7780
rect -1094 7746 -1060 7780
rect -1022 7746 -988 7780
rect -950 7746 -916 7780
rect -878 7746 -844 7780
rect -806 7746 -772 7780
rect -734 7746 -700 7780
rect -662 7746 -628 7780
rect -590 7746 -556 7780
rect -518 7746 -484 7780
rect -446 7746 -412 7780
rect -374 7746 -340 7780
rect -302 7746 -268 7780
rect -230 7746 -196 7780
rect -158 7746 -124 7780
rect -86 7746 -52 7780
rect -14 7746 20 7780
rect 58 7746 92 7780
rect 130 7746 164 7780
rect 202 7746 236 7780
rect 274 7746 308 7780
rect 346 7746 380 7780
rect 418 7746 452 7780
rect 490 7746 524 7780
rect 562 7746 596 7780
rect 634 7746 668 7780
rect 706 7746 740 7780
rect 778 7746 812 7780
rect 850 7746 884 7780
rect 922 7746 956 7780
rect 994 7746 1028 7780
rect 1066 7746 1100 7780
rect 1138 7746 1172 7780
rect 1210 7746 1244 7780
rect 1282 7746 1316 7780
rect 1354 7746 1388 7780
rect 1426 7746 1460 7780
rect 1498 7746 1532 7780
rect 1570 7746 1604 7780
rect -1556 7627 -1522 7661
rect -1556 7555 -1522 7589
rect -1556 7483 -1522 7517
rect -1556 7411 -1522 7445
rect -1556 7339 -1522 7373
rect -1556 7267 -1522 7301
rect -1556 7195 -1522 7229
rect -1556 7123 -1522 7157
rect -1556 7051 -1522 7085
rect 1672 7627 1706 7661
rect 1672 7555 1706 7589
rect 1672 7483 1706 7517
rect 1672 7411 1706 7445
rect 1672 7339 1706 7373
rect 1672 7267 1706 7301
rect 1672 7195 1706 7229
rect 1672 7123 1706 7157
rect 1672 7051 1706 7085
rect -1556 6979 -1522 7013
rect -1556 6907 -1522 6941
rect -1556 6835 -1522 6869
rect -1556 6763 -1522 6797
rect -1556 6691 -1522 6725
rect -1556 6619 -1522 6653
rect -1556 6547 -1522 6581
rect -1556 6475 -1522 6509
rect -1556 6403 -1522 6437
rect -1556 6331 -1522 6365
rect -1556 6259 -1522 6293
rect -1556 6187 -1522 6221
rect -1556 6115 -1522 6149
rect -1556 6043 -1522 6077
rect -1556 5971 -1522 6005
rect -1556 5899 -1522 5933
rect -1556 5827 -1522 5861
rect -1556 5755 -1522 5789
rect -1556 5683 -1522 5717
rect -1556 5611 -1522 5645
rect -1556 5539 -1522 5573
rect -1556 5467 -1522 5501
rect -1556 5395 -1522 5429
rect -1556 5323 -1522 5357
rect -1556 5251 -1522 5285
rect -1556 5179 -1522 5213
rect -1556 5107 -1522 5141
rect -1556 5035 -1522 5069
rect -1556 4963 -1522 4997
rect -1556 4891 -1522 4925
rect -1556 4819 -1522 4853
rect -1556 4747 -1522 4781
rect -1556 4675 -1522 4709
rect -1556 4603 -1522 4637
rect -1556 4531 -1522 4565
rect -1556 4459 -1522 4493
rect -1556 4387 -1522 4421
rect -1556 4315 -1522 4349
rect -1556 4243 -1522 4277
rect -1556 4171 -1522 4205
rect -1556 4099 -1522 4133
rect -1556 4027 -1522 4061
rect -1556 3955 -1522 3989
rect -1556 3883 -1522 3917
rect -1556 3811 -1522 3845
rect -1556 3739 -1522 3773
rect -1556 3667 -1522 3701
rect -1556 3595 -1522 3629
rect -1556 3523 -1522 3557
rect -1556 3451 -1522 3485
rect -1556 3379 -1522 3413
rect -1556 3307 -1522 3341
rect -1556 3235 -1522 3269
rect -1556 3163 -1522 3197
rect -1556 3091 -1522 3125
rect -1556 3019 -1522 3053
rect -1556 2947 -1522 2981
rect -1556 2875 -1522 2909
rect -1556 2803 -1522 2837
rect -1556 2731 -1522 2765
rect -1556 2659 -1522 2693
rect -1556 2587 -1522 2621
rect -1556 2515 -1522 2549
rect -1556 2443 -1522 2477
rect -1556 2371 -1522 2405
rect -1556 2299 -1522 2333
rect -1556 2227 -1522 2261
rect -1556 2155 -1522 2189
rect -1556 2083 -1522 2117
rect -1556 2011 -1522 2045
rect -1556 1939 -1522 1973
rect -1556 1867 -1522 1901
rect -1556 1795 -1522 1829
rect -1556 1723 -1522 1757
rect -1556 1651 -1522 1685
rect -1556 1579 -1522 1613
rect -1556 1507 -1522 1541
rect -1556 1435 -1522 1469
rect -1556 1363 -1522 1397
rect -1556 1291 -1522 1325
rect -1556 1219 -1522 1253
rect -1556 1147 -1522 1181
rect -1556 1075 -1522 1109
rect -1556 1003 -1522 1037
rect -1556 931 -1522 965
rect -1556 859 -1522 893
rect -1556 787 -1522 821
rect -1556 715 -1522 749
rect -1556 643 -1522 677
rect -1556 571 -1522 605
rect -1556 499 -1522 533
rect -1556 427 -1522 461
rect -1556 355 -1522 389
rect -1556 283 -1522 317
rect -1556 211 -1522 245
rect -1556 139 -1522 173
rect -1556 67 -1522 101
rect -1556 -5 -1522 29
rect -1556 -77 -1522 -43
rect -1556 -149 -1522 -115
rect -1556 -221 -1522 -187
rect -1556 -293 -1522 -259
rect -1556 -365 -1522 -331
rect -1556 -437 -1522 -403
rect -1556 -509 -1522 -475
rect -1556 -581 -1522 -547
rect -1556 -653 -1522 -619
rect -1556 -725 -1522 -691
rect -1556 -797 -1522 -763
rect -1556 -869 -1522 -835
rect -1556 -941 -1522 -907
rect -1556 -1013 -1522 -979
rect -554 6820 704 6998
rect -774 6616 -740 6650
rect -774 6544 -740 6578
rect -774 6472 -740 6506
rect -774 6400 -740 6434
rect -774 6328 -740 6362
rect -774 6256 -740 6290
rect -774 6184 -740 6218
rect 890 6616 924 6650
rect 890 6544 924 6578
rect 890 6472 924 6506
rect 890 6400 924 6434
rect 890 6328 924 6362
rect 890 6256 924 6290
rect 890 6184 924 6218
rect -774 6112 -740 6146
rect -774 6040 -740 6074
rect -774 5968 -740 6002
rect -774 5896 -740 5930
rect -774 5824 -740 5858
rect -774 5752 -740 5786
rect -774 5680 -740 5714
rect -774 5608 -740 5642
rect -774 5536 -740 5570
rect -774 5464 -740 5498
rect -774 5392 -740 5426
rect -774 5320 -740 5354
rect -774 5248 -740 5282
rect -774 5176 -740 5210
rect -774 5104 -740 5138
rect -774 5032 -740 5066
rect -774 4960 -740 4994
rect -774 4888 -740 4922
rect -774 4816 -740 4850
rect -774 4744 -740 4778
rect -774 4672 -740 4706
rect -774 4600 -740 4634
rect -774 4528 -740 4562
rect -774 4456 -740 4490
rect -774 4384 -740 4418
rect -774 4312 -740 4346
rect -774 4240 -740 4274
rect -774 4168 -740 4202
rect -774 4096 -740 4130
rect -774 4024 -740 4058
rect -774 3952 -740 3986
rect -774 3880 -740 3914
rect -774 3808 -740 3842
rect -774 3736 -740 3770
rect -774 3664 -740 3698
rect -774 3592 -740 3626
rect -774 3520 -740 3554
rect -774 3448 -740 3482
rect -774 3376 -740 3410
rect -774 3304 -740 3338
rect -774 3232 -740 3266
rect -774 3160 -740 3194
rect -774 3088 -740 3122
rect -774 3016 -740 3050
rect -774 2944 -740 2978
rect -774 2872 -740 2906
rect -774 2800 -740 2834
rect -774 2728 -740 2762
rect -774 2656 -740 2690
rect -774 2584 -740 2618
rect -774 2512 -740 2546
rect -774 2440 -740 2474
rect -774 2368 -740 2402
rect -774 2296 -740 2330
rect -774 2224 -740 2258
rect -774 2152 -740 2186
rect -774 2080 -740 2114
rect -774 2008 -740 2042
rect -774 1936 -740 1970
rect -774 1864 -740 1898
rect -774 1792 -740 1826
rect -774 1720 -740 1754
rect -774 1648 -740 1682
rect -774 1576 -740 1610
rect -774 1504 -740 1538
rect -774 1432 -740 1466
rect -774 1360 -740 1394
rect -774 1288 -740 1322
rect -774 1216 -740 1250
rect -774 1144 -740 1178
rect -774 1072 -740 1106
rect -774 1000 -740 1034
rect -774 928 -740 962
rect -774 856 -740 890
rect -774 784 -740 818
rect -774 712 -740 746
rect -774 640 -740 674
rect -774 568 -740 602
rect -774 496 -740 530
rect -774 424 -740 458
rect -774 352 -740 386
rect -774 280 -740 314
rect -774 208 -740 242
rect -774 136 -740 170
rect -774 64 -740 98
rect -774 -8 -740 26
rect -774 -80 -740 -46
rect -774 -152 -740 -118
rect -647 -152 -469 6146
rect -122 -152 272 6146
rect 619 -152 797 6146
rect 890 6112 924 6146
rect 890 6040 924 6074
rect 890 5968 924 6002
rect 890 5896 924 5930
rect 890 5824 924 5858
rect 890 5752 924 5786
rect 890 5680 924 5714
rect 890 5608 924 5642
rect 890 5536 924 5570
rect 890 5464 924 5498
rect 890 5392 924 5426
rect 890 5320 924 5354
rect 890 5248 924 5282
rect 890 5176 924 5210
rect 890 5104 924 5138
rect 890 5032 924 5066
rect 890 4960 924 4994
rect 890 4888 924 4922
rect 890 4816 924 4850
rect 890 4744 924 4778
rect 890 4672 924 4706
rect 890 4600 924 4634
rect 890 4528 924 4562
rect 890 4456 924 4490
rect 890 4384 924 4418
rect 890 4312 924 4346
rect 890 4240 924 4274
rect 890 4168 924 4202
rect 890 4096 924 4130
rect 890 4024 924 4058
rect 890 3952 924 3986
rect 890 3880 924 3914
rect 890 3808 924 3842
rect 890 3736 924 3770
rect 890 3664 924 3698
rect 890 3592 924 3626
rect 890 3520 924 3554
rect 890 3448 924 3482
rect 890 3376 924 3410
rect 890 3304 924 3338
rect 890 3232 924 3266
rect 890 3160 924 3194
rect 890 3088 924 3122
rect 890 3016 924 3050
rect 890 2944 924 2978
rect 890 2872 924 2906
rect 890 2800 924 2834
rect 890 2728 924 2762
rect 890 2656 924 2690
rect 890 2584 924 2618
rect 890 2512 924 2546
rect 890 2440 924 2474
rect 890 2368 924 2402
rect 890 2296 924 2330
rect 890 2224 924 2258
rect 890 2152 924 2186
rect 890 2080 924 2114
rect 890 2008 924 2042
rect 890 1936 924 1970
rect 890 1864 924 1898
rect 890 1792 924 1826
rect 890 1720 924 1754
rect 890 1648 924 1682
rect 890 1576 924 1610
rect 890 1504 924 1538
rect 890 1432 924 1466
rect 890 1360 924 1394
rect 890 1288 924 1322
rect 890 1216 924 1250
rect 890 1144 924 1178
rect 890 1072 924 1106
rect 890 1000 924 1034
rect 890 928 924 962
rect 890 856 924 890
rect 890 784 924 818
rect 890 712 924 746
rect 890 640 924 674
rect 890 568 924 602
rect 890 496 924 530
rect 890 424 924 458
rect 890 352 924 386
rect 890 280 924 314
rect 890 208 924 242
rect 890 136 924 170
rect 890 64 924 98
rect 890 -8 924 26
rect 890 -80 924 -46
rect 890 -152 924 -118
rect -774 -224 -740 -190
rect -774 -296 -740 -262
rect -774 -368 -740 -334
rect -774 -440 -740 -406
rect 890 -224 924 -190
rect 890 -296 924 -262
rect 890 -368 924 -334
rect 890 -440 924 -406
rect -774 -512 -740 -478
rect -774 -584 -740 -550
rect -774 -656 -740 -622
rect -130 -493 -96 -459
rect -56 -493 -22 -459
rect 18 -493 52 -459
rect 92 -493 126 -459
rect 166 -493 200 -459
rect 240 -493 274 -459
rect -130 -567 -96 -533
rect -56 -567 -22 -533
rect 18 -567 52 -533
rect 92 -567 126 -533
rect 166 -567 200 -533
rect 240 -567 274 -533
rect -130 -641 -96 -607
rect -56 -641 -22 -607
rect 18 -641 52 -607
rect 92 -641 126 -607
rect 166 -641 200 -607
rect 240 -641 274 -607
rect 890 -512 924 -478
rect 890 -584 924 -550
rect 890 -656 924 -622
rect -554 -998 704 -820
rect 1672 6979 1706 7013
rect 1672 6907 1706 6941
rect 1672 6835 1706 6869
rect 1672 6763 1706 6797
rect 1672 6691 1706 6725
rect 1672 6619 1706 6653
rect 1672 6547 1706 6581
rect 1672 6475 1706 6509
rect 1672 6403 1706 6437
rect 1672 6331 1706 6365
rect 1672 6259 1706 6293
rect 1672 6187 1706 6221
rect 1672 6115 1706 6149
rect 1672 6043 1706 6077
rect 1672 5971 1706 6005
rect 1672 5899 1706 5933
rect 1672 5827 1706 5861
rect 1672 5755 1706 5789
rect 1672 5683 1706 5717
rect 1672 5611 1706 5645
rect 1672 5539 1706 5573
rect 1672 5467 1706 5501
rect 1672 5395 1706 5429
rect 1672 5323 1706 5357
rect 1672 5251 1706 5285
rect 1672 5179 1706 5213
rect 1672 5107 1706 5141
rect 1672 5035 1706 5069
rect 1672 4963 1706 4997
rect 1672 4891 1706 4925
rect 1672 4819 1706 4853
rect 1672 4747 1706 4781
rect 1672 4675 1706 4709
rect 1672 4603 1706 4637
rect 1672 4531 1706 4565
rect 1672 4459 1706 4493
rect 1672 4387 1706 4421
rect 1672 4315 1706 4349
rect 1672 4243 1706 4277
rect 1672 4171 1706 4205
rect 1672 4099 1706 4133
rect 1672 4027 1706 4061
rect 1672 3955 1706 3989
rect 1672 3883 1706 3917
rect 1672 3811 1706 3845
rect 1672 3739 1706 3773
rect 1672 3667 1706 3701
rect 1672 3595 1706 3629
rect 1672 3523 1706 3557
rect 1672 3451 1706 3485
rect 1672 3379 1706 3413
rect 1672 3307 1706 3341
rect 1672 3235 1706 3269
rect 1672 3163 1706 3197
rect 1672 3091 1706 3125
rect 1672 3019 1706 3053
rect 1672 2947 1706 2981
rect 1672 2875 1706 2909
rect 1672 2803 1706 2837
rect 1672 2731 1706 2765
rect 1672 2659 1706 2693
rect 1672 2587 1706 2621
rect 1672 2515 1706 2549
rect 1672 2443 1706 2477
rect 1672 2371 1706 2405
rect 1672 2299 1706 2333
rect 1672 2227 1706 2261
rect 1672 2155 1706 2189
rect 1672 2083 1706 2117
rect 1672 2011 1706 2045
rect 1672 1939 1706 1973
rect 1672 1867 1706 1901
rect 1672 1795 1706 1829
rect 1672 1723 1706 1757
rect 1672 1651 1706 1685
rect 1672 1579 1706 1613
rect 1672 1507 1706 1541
rect 1672 1435 1706 1469
rect 1672 1363 1706 1397
rect 1672 1291 1706 1325
rect 1672 1219 1706 1253
rect 1672 1147 1706 1181
rect 1672 1075 1706 1109
rect 1672 1003 1706 1037
rect 1672 931 1706 965
rect 1672 859 1706 893
rect 1672 787 1706 821
rect 1672 715 1706 749
rect 1672 643 1706 677
rect 1672 571 1706 605
rect 1672 499 1706 533
rect 1672 427 1706 461
rect 1672 355 1706 389
rect 1672 283 1706 317
rect 1672 211 1706 245
rect 1672 139 1706 173
rect 1672 67 1706 101
rect 1672 -5 1706 29
rect 1672 -77 1706 -43
rect 1672 -149 1706 -115
rect 1672 -221 1706 -187
rect 1672 -293 1706 -259
rect 1672 -365 1706 -331
rect 1672 -437 1706 -403
rect 1672 -509 1706 -475
rect 1672 -581 1706 -547
rect 1672 -653 1706 -619
rect 1672 -725 1706 -691
rect 1672 -797 1706 -763
rect 1672 -869 1706 -835
rect 1672 -941 1706 -907
rect 1672 -1013 1706 -979
rect -1556 -1085 -1522 -1051
rect -1556 -1157 -1522 -1123
rect -1556 -1229 -1522 -1195
rect -1556 -1301 -1522 -1267
rect -1556 -1373 -1522 -1339
rect -1556 -1445 -1522 -1411
rect -1556 -1517 -1522 -1483
rect -1556 -1589 -1522 -1555
rect -1556 -1661 -1522 -1627
rect 1672 -1085 1706 -1051
rect 1672 -1157 1706 -1123
rect 1672 -1229 1706 -1195
rect 1672 -1301 1706 -1267
rect 1672 -1373 1706 -1339
rect 1672 -1445 1706 -1411
rect 1672 -1517 1706 -1483
rect 1672 -1589 1706 -1555
rect 1672 -1661 1706 -1627
rect -1454 -1780 -1420 -1746
rect -1382 -1780 -1348 -1746
rect -1310 -1780 -1276 -1746
rect -1238 -1780 -1204 -1746
rect -1166 -1780 -1132 -1746
rect -1094 -1780 -1060 -1746
rect -1022 -1780 -988 -1746
rect -950 -1780 -916 -1746
rect -878 -1780 -844 -1746
rect -806 -1780 -772 -1746
rect -734 -1780 -700 -1746
rect -662 -1780 -628 -1746
rect -590 -1780 -556 -1746
rect -518 -1780 -484 -1746
rect -446 -1780 -412 -1746
rect -374 -1780 -340 -1746
rect -302 -1780 -268 -1746
rect -230 -1780 -196 -1746
rect -158 -1780 -124 -1746
rect -86 -1780 -52 -1746
rect -14 -1780 20 -1746
rect 58 -1780 92 -1746
rect 130 -1780 164 -1746
rect 202 -1780 236 -1746
rect 274 -1780 308 -1746
rect 346 -1780 380 -1746
rect 418 -1780 452 -1746
rect 490 -1780 524 -1746
rect 562 -1780 596 -1746
rect 634 -1780 668 -1746
rect 706 -1780 740 -1746
rect 778 -1780 812 -1746
rect 850 -1780 884 -1746
rect 922 -1780 956 -1746
rect 994 -1780 1028 -1746
rect 1066 -1780 1100 -1746
rect 1138 -1780 1172 -1746
rect 1210 -1780 1244 -1746
rect 1282 -1780 1316 -1746
rect 1354 -1780 1388 -1746
rect 1426 -1780 1460 -1746
rect 1498 -1780 1532 -1746
rect 1570 -1780 1604 -1746
<< metal1 >>
rect -1580 7780 1730 7804
rect -1580 7746 -1454 7780
rect -1420 7746 -1382 7780
rect -1348 7746 -1310 7780
rect -1276 7746 -1238 7780
rect -1204 7746 -1166 7780
rect -1132 7746 -1094 7780
rect -1060 7746 -1022 7780
rect -988 7746 -950 7780
rect -916 7746 -878 7780
rect -844 7746 -806 7780
rect -772 7746 -734 7780
rect -700 7746 -662 7780
rect -628 7746 -590 7780
rect -556 7746 -518 7780
rect -484 7746 -446 7780
rect -412 7746 -374 7780
rect -340 7746 -302 7780
rect -268 7746 -230 7780
rect -196 7746 -158 7780
rect -124 7746 -86 7780
rect -52 7746 -14 7780
rect 20 7746 58 7780
rect 92 7746 130 7780
rect 164 7746 202 7780
rect 236 7746 274 7780
rect 308 7746 346 7780
rect 380 7746 418 7780
rect 452 7746 490 7780
rect 524 7746 562 7780
rect 596 7746 634 7780
rect 668 7746 706 7780
rect 740 7746 778 7780
rect 812 7746 850 7780
rect 884 7746 922 7780
rect 956 7746 994 7780
rect 1028 7746 1066 7780
rect 1100 7746 1138 7780
rect 1172 7746 1210 7780
rect 1244 7746 1282 7780
rect 1316 7746 1354 7780
rect 1388 7746 1426 7780
rect 1460 7746 1498 7780
rect 1532 7746 1570 7780
rect 1604 7746 1730 7780
rect -1580 7722 1730 7746
rect -1580 7661 -1498 7722
rect -1580 7627 -1556 7661
rect -1522 7627 -1498 7661
rect -1580 7589 -1498 7627
rect -1580 7555 -1556 7589
rect -1522 7555 -1498 7589
rect -1580 7517 -1498 7555
rect -1580 7483 -1556 7517
rect -1522 7483 -1498 7517
rect -1580 7445 -1498 7483
rect -1580 7411 -1556 7445
rect -1522 7411 -1498 7445
rect -1580 7373 -1498 7411
rect -1580 7339 -1556 7373
rect -1522 7339 -1498 7373
rect -1580 7301 -1498 7339
rect -1580 7267 -1556 7301
rect -1522 7267 -1498 7301
rect -1580 7229 -1498 7267
rect -1580 7195 -1556 7229
rect -1522 7195 -1498 7229
rect -1580 7157 -1498 7195
rect -1580 7123 -1556 7157
rect -1522 7123 -1498 7157
rect -1580 7085 -1498 7123
rect -1580 7051 -1556 7085
rect -1522 7051 -1498 7085
rect -1580 7013 -1498 7051
rect 1648 7661 1730 7722
rect 1648 7627 1672 7661
rect 1706 7627 1730 7661
rect 1648 7589 1730 7627
rect 1648 7555 1672 7589
rect 1706 7555 1730 7589
rect 1648 7517 1730 7555
rect 1648 7483 1672 7517
rect 1706 7483 1730 7517
rect 1648 7445 1730 7483
rect 1648 7411 1672 7445
rect 1706 7411 1730 7445
rect 1648 7373 1730 7411
rect 1648 7339 1672 7373
rect 1706 7339 1730 7373
rect 1648 7301 1730 7339
rect 1648 7267 1672 7301
rect 1706 7267 1730 7301
rect 1648 7229 1730 7267
rect 1648 7195 1672 7229
rect 1706 7195 1730 7229
rect 1648 7157 1730 7195
rect 1648 7123 1672 7157
rect 1706 7123 1730 7157
rect 1648 7085 1730 7123
rect 1648 7051 1672 7085
rect 1706 7051 1730 7085
rect -1580 6979 -1556 7013
rect -1522 6979 -1498 7013
rect -1580 6941 -1498 6979
rect -1580 6907 -1556 6941
rect -1522 6907 -1498 6941
rect -1580 6869 -1498 6907
rect -1580 6835 -1556 6869
rect -1522 6835 -1498 6869
rect -1580 6797 -1498 6835
rect -1580 6763 -1556 6797
rect -1522 6763 -1498 6797
rect -1580 6725 -1498 6763
rect -1580 6691 -1556 6725
rect -1522 6691 -1498 6725
rect -1580 6653 -1498 6691
rect -1580 6619 -1556 6653
rect -1522 6619 -1498 6653
rect -1580 6581 -1498 6619
rect -1580 6547 -1556 6581
rect -1522 6547 -1498 6581
rect -1580 6509 -1498 6547
rect -1580 6475 -1556 6509
rect -1522 6475 -1498 6509
rect -1580 6437 -1498 6475
rect -1580 6403 -1556 6437
rect -1522 6403 -1498 6437
rect -1580 6365 -1498 6403
rect -1580 6331 -1556 6365
rect -1522 6331 -1498 6365
rect -1580 6293 -1498 6331
rect -1580 6259 -1556 6293
rect -1522 6259 -1498 6293
rect -1580 6221 -1498 6259
rect -1580 6187 -1556 6221
rect -1522 6187 -1498 6221
rect -1580 6149 -1498 6187
rect -1580 6115 -1556 6149
rect -1522 6115 -1498 6149
rect -1580 6077 -1498 6115
rect -1580 6043 -1556 6077
rect -1522 6043 -1498 6077
rect -1580 6005 -1498 6043
rect -1580 5971 -1556 6005
rect -1522 5971 -1498 6005
rect -1580 5933 -1498 5971
rect -1580 5899 -1556 5933
rect -1522 5899 -1498 5933
rect -1580 5861 -1498 5899
rect -1580 5827 -1556 5861
rect -1522 5827 -1498 5861
rect -1580 5789 -1498 5827
rect -1580 5755 -1556 5789
rect -1522 5755 -1498 5789
rect -1580 5717 -1498 5755
rect -1580 5683 -1556 5717
rect -1522 5683 -1498 5717
rect -1580 5645 -1498 5683
rect -1580 5611 -1556 5645
rect -1522 5611 -1498 5645
rect -1580 5573 -1498 5611
rect -1580 5539 -1556 5573
rect -1522 5539 -1498 5573
rect -1580 5501 -1498 5539
rect -1580 5467 -1556 5501
rect -1522 5467 -1498 5501
rect -1580 5429 -1498 5467
rect -1580 5395 -1556 5429
rect -1522 5395 -1498 5429
rect -1580 5357 -1498 5395
rect -1580 5323 -1556 5357
rect -1522 5323 -1498 5357
rect -1580 5285 -1498 5323
rect -1580 5251 -1556 5285
rect -1522 5251 -1498 5285
rect -1580 5213 -1498 5251
rect -1580 5179 -1556 5213
rect -1522 5179 -1498 5213
rect -1580 5141 -1498 5179
rect -1580 5107 -1556 5141
rect -1522 5107 -1498 5141
rect -1580 5069 -1498 5107
rect -1580 5035 -1556 5069
rect -1522 5035 -1498 5069
rect -1580 4997 -1498 5035
rect -1580 4963 -1556 4997
rect -1522 4963 -1498 4997
rect -1580 4925 -1498 4963
rect -1580 4891 -1556 4925
rect -1522 4891 -1498 4925
rect -1580 4853 -1498 4891
rect -1580 4819 -1556 4853
rect -1522 4819 -1498 4853
rect -1580 4781 -1498 4819
rect -1580 4747 -1556 4781
rect -1522 4747 -1498 4781
rect -1580 4709 -1498 4747
rect -1580 4675 -1556 4709
rect -1522 4675 -1498 4709
rect -1580 4637 -1498 4675
rect -1580 4603 -1556 4637
rect -1522 4603 -1498 4637
rect -1580 4565 -1498 4603
rect -1580 4531 -1556 4565
rect -1522 4531 -1498 4565
rect -1580 4493 -1498 4531
rect -1580 4459 -1556 4493
rect -1522 4459 -1498 4493
rect -1580 4421 -1498 4459
rect -1580 4387 -1556 4421
rect -1522 4387 -1498 4421
rect -1580 4349 -1498 4387
rect -1580 4315 -1556 4349
rect -1522 4315 -1498 4349
rect -1580 4277 -1498 4315
rect -1580 4243 -1556 4277
rect -1522 4243 -1498 4277
rect -1580 4205 -1498 4243
rect -1580 4171 -1556 4205
rect -1522 4171 -1498 4205
rect -1580 4133 -1498 4171
rect -1580 4099 -1556 4133
rect -1522 4099 -1498 4133
rect -1580 4061 -1498 4099
rect -1580 4027 -1556 4061
rect -1522 4027 -1498 4061
rect -1580 3989 -1498 4027
rect -1580 3955 -1556 3989
rect -1522 3955 -1498 3989
rect -1580 3917 -1498 3955
rect -1580 3883 -1556 3917
rect -1522 3883 -1498 3917
rect -1580 3845 -1498 3883
rect -1580 3811 -1556 3845
rect -1522 3811 -1498 3845
rect -1580 3773 -1498 3811
rect -1580 3739 -1556 3773
rect -1522 3739 -1498 3773
rect -1580 3701 -1498 3739
rect -1580 3667 -1556 3701
rect -1522 3667 -1498 3701
rect -1580 3629 -1498 3667
rect -1580 3595 -1556 3629
rect -1522 3595 -1498 3629
rect -1580 3557 -1498 3595
rect -1580 3523 -1556 3557
rect -1522 3523 -1498 3557
rect -1580 3485 -1498 3523
rect -1580 3451 -1556 3485
rect -1522 3451 -1498 3485
rect -1580 3413 -1498 3451
rect -1580 3379 -1556 3413
rect -1522 3379 -1498 3413
rect -1580 3341 -1498 3379
rect -1580 3307 -1556 3341
rect -1522 3307 -1498 3341
rect -1580 3269 -1498 3307
rect -1580 3235 -1556 3269
rect -1522 3235 -1498 3269
rect -1580 3197 -1498 3235
rect -1580 3163 -1556 3197
rect -1522 3163 -1498 3197
rect -1580 3125 -1498 3163
rect -1580 3091 -1556 3125
rect -1522 3091 -1498 3125
rect -1580 3053 -1498 3091
rect -1580 3019 -1556 3053
rect -1522 3019 -1498 3053
rect -1580 2981 -1498 3019
rect -1580 2947 -1556 2981
rect -1522 2947 -1498 2981
rect -1580 2909 -1498 2947
rect -1580 2875 -1556 2909
rect -1522 2875 -1498 2909
rect -1580 2837 -1498 2875
rect -1580 2803 -1556 2837
rect -1522 2803 -1498 2837
rect -1580 2765 -1498 2803
rect -1580 2731 -1556 2765
rect -1522 2731 -1498 2765
rect -1580 2693 -1498 2731
rect -1580 2659 -1556 2693
rect -1522 2659 -1498 2693
rect -1580 2621 -1498 2659
rect -1580 2587 -1556 2621
rect -1522 2587 -1498 2621
rect -1580 2549 -1498 2587
rect -1580 2515 -1556 2549
rect -1522 2515 -1498 2549
rect -1580 2477 -1498 2515
rect -1580 2443 -1556 2477
rect -1522 2443 -1498 2477
rect -1580 2405 -1498 2443
rect -1580 2371 -1556 2405
rect -1522 2371 -1498 2405
rect -1580 2333 -1498 2371
rect -1580 2299 -1556 2333
rect -1522 2299 -1498 2333
rect -1580 2261 -1498 2299
rect -1580 2227 -1556 2261
rect -1522 2227 -1498 2261
rect -1580 2189 -1498 2227
rect -1580 2155 -1556 2189
rect -1522 2155 -1498 2189
rect -1580 2117 -1498 2155
rect -1580 2083 -1556 2117
rect -1522 2083 -1498 2117
rect -1580 2045 -1498 2083
rect -1580 2011 -1556 2045
rect -1522 2011 -1498 2045
rect -1580 1973 -1498 2011
rect -1580 1939 -1556 1973
rect -1522 1939 -1498 1973
rect -1580 1901 -1498 1939
rect -1580 1867 -1556 1901
rect -1522 1867 -1498 1901
rect -1580 1829 -1498 1867
rect -1580 1795 -1556 1829
rect -1522 1795 -1498 1829
rect -1580 1757 -1498 1795
rect -1580 1723 -1556 1757
rect -1522 1723 -1498 1757
rect -1580 1685 -1498 1723
rect -1580 1651 -1556 1685
rect -1522 1651 -1498 1685
rect -1580 1613 -1498 1651
rect -1580 1579 -1556 1613
rect -1522 1579 -1498 1613
rect -1580 1541 -1498 1579
rect -1580 1507 -1556 1541
rect -1522 1507 -1498 1541
rect -1580 1469 -1498 1507
rect -1580 1435 -1556 1469
rect -1522 1435 -1498 1469
rect -1580 1397 -1498 1435
rect -1580 1363 -1556 1397
rect -1522 1363 -1498 1397
rect -1580 1325 -1498 1363
rect -1580 1291 -1556 1325
rect -1522 1291 -1498 1325
rect -1580 1253 -1498 1291
rect -1580 1219 -1556 1253
rect -1522 1219 -1498 1253
rect -1580 1181 -1498 1219
rect -1580 1147 -1556 1181
rect -1522 1147 -1498 1181
rect -1580 1109 -1498 1147
rect -1580 1075 -1556 1109
rect -1522 1075 -1498 1109
rect -1580 1037 -1498 1075
rect -1580 1003 -1556 1037
rect -1522 1003 -1498 1037
rect -1580 965 -1498 1003
rect -1580 931 -1556 965
rect -1522 931 -1498 965
rect -1580 893 -1498 931
rect -1580 859 -1556 893
rect -1522 859 -1498 893
rect -1580 821 -1498 859
rect -1580 787 -1556 821
rect -1522 787 -1498 821
rect -1580 749 -1498 787
rect -1580 715 -1556 749
rect -1522 715 -1498 749
rect -1580 677 -1498 715
rect -1580 643 -1556 677
rect -1522 643 -1498 677
rect -1580 605 -1498 643
rect -1580 571 -1556 605
rect -1522 571 -1498 605
rect -1580 533 -1498 571
rect -1580 499 -1556 533
rect -1522 499 -1498 533
rect -1580 461 -1498 499
rect -1580 427 -1556 461
rect -1522 427 -1498 461
rect -1580 389 -1498 427
rect -1580 355 -1556 389
rect -1522 355 -1498 389
rect -1580 317 -1498 355
rect -1580 283 -1556 317
rect -1522 283 -1498 317
rect -1580 245 -1498 283
rect -1580 211 -1556 245
rect -1522 211 -1498 245
rect -1580 173 -1498 211
rect -1580 139 -1556 173
rect -1522 139 -1498 173
rect -1580 101 -1498 139
rect -1580 67 -1556 101
rect -1522 67 -1498 101
rect -1580 29 -1498 67
rect -1580 -5 -1556 29
rect -1522 -5 -1498 29
rect -1580 -43 -1498 -5
rect -1580 -77 -1556 -43
rect -1522 -77 -1498 -43
rect -1580 -115 -1498 -77
rect -1580 -149 -1556 -115
rect -1522 -149 -1498 -115
rect -1580 -187 -1498 -149
rect -1580 -221 -1556 -187
rect -1522 -221 -1498 -187
rect -1580 -259 -1498 -221
rect -1580 -293 -1556 -259
rect -1522 -293 -1498 -259
rect -1580 -331 -1498 -293
rect -1580 -365 -1556 -331
rect -1522 -365 -1498 -331
rect -1580 -403 -1498 -365
rect -1580 -437 -1556 -403
rect -1522 -437 -1498 -403
rect -1580 -475 -1498 -437
rect -1580 -509 -1556 -475
rect -1522 -509 -1498 -475
rect -1580 -547 -1498 -509
rect -1580 -581 -1556 -547
rect -1522 -581 -1498 -547
rect -1580 -619 -1498 -581
rect -1580 -653 -1556 -619
rect -1522 -653 -1498 -619
rect -1580 -691 -1498 -653
rect -1580 -725 -1556 -691
rect -1522 -725 -1498 -691
rect -1580 -763 -1498 -725
rect -1580 -797 -1556 -763
rect -1522 -797 -1498 -763
rect -1580 -835 -1498 -797
rect -1580 -869 -1556 -835
rect -1522 -869 -1498 -835
rect -1580 -907 -1498 -869
rect -1580 -941 -1556 -907
rect -1522 -941 -1498 -907
rect -1580 -979 -1498 -941
rect -1580 -1013 -1556 -979
rect -1522 -1013 -1498 -979
rect -1580 -1051 -1498 -1013
rect -798 6998 948 7022
rect -798 6820 -554 6998
rect 704 6820 948 6998
rect -798 6757 948 6820
rect -798 6650 -716 6757
rect -798 6616 -774 6650
rect -740 6616 -716 6650
rect -798 6578 -716 6616
rect -798 6544 -774 6578
rect -740 6544 -716 6578
rect -798 6506 -716 6544
rect -798 6472 -774 6506
rect -740 6472 -716 6506
rect -798 6434 -716 6472
rect -798 6400 -774 6434
rect -740 6400 -716 6434
rect -798 6362 -716 6400
rect -798 6328 -774 6362
rect -740 6328 -716 6362
rect -798 6290 -716 6328
rect -798 6256 -774 6290
rect -740 6256 -716 6290
rect -798 6218 -716 6256
rect -798 6184 -774 6218
rect -740 6184 -716 6218
rect -798 6146 -716 6184
rect 866 6650 948 6757
rect 866 6616 890 6650
rect 924 6616 948 6650
rect 866 6578 948 6616
rect 866 6544 890 6578
rect 924 6544 948 6578
rect 866 6506 948 6544
rect 866 6472 890 6506
rect 924 6472 948 6506
rect 866 6434 948 6472
rect 866 6400 890 6434
rect 924 6400 948 6434
rect 866 6362 948 6400
rect 866 6328 890 6362
rect 924 6328 948 6362
rect 866 6290 948 6328
rect 866 6256 890 6290
rect 924 6256 948 6290
rect 866 6218 948 6256
rect 866 6184 890 6218
rect 924 6184 948 6218
rect -798 6112 -774 6146
rect -740 6112 -716 6146
rect -798 6074 -716 6112
rect -798 6040 -774 6074
rect -740 6040 -716 6074
rect -798 6002 -716 6040
rect -798 5968 -774 6002
rect -740 5968 -716 6002
rect -798 5930 -716 5968
rect -798 5896 -774 5930
rect -740 5896 -716 5930
rect -798 5858 -716 5896
rect -798 5824 -774 5858
rect -740 5824 -716 5858
rect -798 5786 -716 5824
rect -798 5752 -774 5786
rect -740 5752 -716 5786
rect -798 5714 -716 5752
rect -798 5680 -774 5714
rect -740 5680 -716 5714
rect -798 5642 -716 5680
rect -798 5608 -774 5642
rect -740 5608 -716 5642
rect -798 5570 -716 5608
rect -798 5536 -774 5570
rect -740 5536 -716 5570
rect -798 5498 -716 5536
rect -798 5464 -774 5498
rect -740 5464 -716 5498
rect -798 5426 -716 5464
rect -798 5392 -774 5426
rect -740 5392 -716 5426
rect -798 5354 -716 5392
rect -798 5320 -774 5354
rect -740 5320 -716 5354
rect -798 5282 -716 5320
rect -798 5248 -774 5282
rect -740 5248 -716 5282
rect -798 5210 -716 5248
rect -798 5176 -774 5210
rect -740 5176 -716 5210
rect -798 5138 -716 5176
rect -798 5104 -774 5138
rect -740 5104 -716 5138
rect -798 5066 -716 5104
rect -798 5032 -774 5066
rect -740 5032 -716 5066
rect -798 4994 -716 5032
rect -798 4960 -774 4994
rect -740 4960 -716 4994
rect -798 4922 -716 4960
rect -798 4888 -774 4922
rect -740 4888 -716 4922
rect -798 4850 -716 4888
rect -798 4816 -774 4850
rect -740 4816 -716 4850
rect -798 4778 -716 4816
rect -798 4744 -774 4778
rect -740 4744 -716 4778
rect -798 4706 -716 4744
rect -798 4672 -774 4706
rect -740 4672 -716 4706
rect -798 4634 -716 4672
rect -798 4600 -774 4634
rect -740 4600 -716 4634
rect -798 4562 -716 4600
rect -798 4528 -774 4562
rect -740 4528 -716 4562
rect -798 4490 -716 4528
rect -798 4456 -774 4490
rect -740 4456 -716 4490
rect -798 4418 -716 4456
rect -798 4384 -774 4418
rect -740 4384 -716 4418
rect -798 4346 -716 4384
rect -798 4312 -774 4346
rect -740 4312 -716 4346
rect -798 4274 -716 4312
rect -798 4240 -774 4274
rect -740 4240 -716 4274
rect -798 4202 -716 4240
rect -798 4168 -774 4202
rect -740 4168 -716 4202
rect -798 4130 -716 4168
rect -798 4096 -774 4130
rect -740 4096 -716 4130
rect -798 4058 -716 4096
rect -798 4024 -774 4058
rect -740 4024 -716 4058
rect -798 3986 -716 4024
rect -798 3952 -774 3986
rect -740 3952 -716 3986
rect -798 3914 -716 3952
rect -798 3880 -774 3914
rect -740 3880 -716 3914
rect -798 3842 -716 3880
rect -798 3808 -774 3842
rect -740 3808 -716 3842
rect -798 3770 -716 3808
rect -798 3736 -774 3770
rect -740 3736 -716 3770
rect -798 3698 -716 3736
rect -798 3664 -774 3698
rect -740 3664 -716 3698
rect -798 3626 -716 3664
rect -798 3592 -774 3626
rect -740 3592 -716 3626
rect -798 3554 -716 3592
rect -798 3520 -774 3554
rect -740 3520 -716 3554
rect -798 3482 -716 3520
rect -798 3448 -774 3482
rect -740 3448 -716 3482
rect -798 3410 -716 3448
rect -798 3376 -774 3410
rect -740 3376 -716 3410
rect -798 3338 -716 3376
rect -798 3304 -774 3338
rect -740 3304 -716 3338
rect -798 3266 -716 3304
rect -798 3232 -774 3266
rect -740 3232 -716 3266
rect -798 3194 -716 3232
rect -798 3160 -774 3194
rect -740 3160 -716 3194
rect -798 3122 -716 3160
rect -798 3088 -774 3122
rect -740 3088 -716 3122
rect -798 3050 -716 3088
rect -798 3016 -774 3050
rect -740 3016 -716 3050
rect -798 2978 -716 3016
rect -798 2944 -774 2978
rect -740 2944 -716 2978
rect -798 2906 -716 2944
rect -798 2872 -774 2906
rect -740 2872 -716 2906
rect -798 2834 -716 2872
rect -798 2800 -774 2834
rect -740 2800 -716 2834
rect -798 2762 -716 2800
rect -798 2728 -774 2762
rect -740 2728 -716 2762
rect -798 2690 -716 2728
rect -798 2656 -774 2690
rect -740 2656 -716 2690
rect -798 2618 -716 2656
rect -798 2584 -774 2618
rect -740 2584 -716 2618
rect -798 2546 -716 2584
rect -798 2512 -774 2546
rect -740 2512 -716 2546
rect -798 2474 -716 2512
rect -798 2440 -774 2474
rect -740 2440 -716 2474
rect -798 2402 -716 2440
rect -798 2368 -774 2402
rect -740 2368 -716 2402
rect -798 2330 -716 2368
rect -798 2296 -774 2330
rect -740 2296 -716 2330
rect -798 2258 -716 2296
rect -798 2224 -774 2258
rect -740 2224 -716 2258
rect -798 2186 -716 2224
rect -798 2152 -774 2186
rect -740 2152 -716 2186
rect -798 2114 -716 2152
rect -798 2080 -774 2114
rect -740 2080 -716 2114
rect -798 2042 -716 2080
rect -798 2008 -774 2042
rect -740 2008 -716 2042
rect -798 1970 -716 2008
rect -798 1936 -774 1970
rect -740 1936 -716 1970
rect -798 1898 -716 1936
rect -798 1864 -774 1898
rect -740 1864 -716 1898
rect -798 1826 -716 1864
rect -798 1792 -774 1826
rect -740 1792 -716 1826
rect -798 1754 -716 1792
rect -798 1720 -774 1754
rect -740 1720 -716 1754
rect -798 1682 -716 1720
rect -798 1648 -774 1682
rect -740 1648 -716 1682
rect -798 1610 -716 1648
rect -798 1576 -774 1610
rect -740 1576 -716 1610
rect -798 1538 -716 1576
rect -798 1504 -774 1538
rect -740 1504 -716 1538
rect -798 1466 -716 1504
rect -798 1432 -774 1466
rect -740 1432 -716 1466
rect -798 1394 -716 1432
rect -798 1360 -774 1394
rect -740 1360 -716 1394
rect -798 1322 -716 1360
rect -798 1288 -774 1322
rect -740 1288 -716 1322
rect -798 1250 -716 1288
rect -798 1216 -774 1250
rect -740 1216 -716 1250
rect -798 1178 -716 1216
rect -798 1144 -774 1178
rect -740 1144 -716 1178
rect -798 1106 -716 1144
rect -798 1072 -774 1106
rect -740 1072 -716 1106
rect -798 1034 -716 1072
rect -798 1000 -774 1034
rect -740 1000 -716 1034
rect -798 962 -716 1000
rect -798 928 -774 962
rect -740 928 -716 962
rect -798 890 -716 928
rect -798 856 -774 890
rect -740 856 -716 890
rect -798 818 -716 856
rect -798 784 -774 818
rect -740 784 -716 818
rect -798 746 -716 784
rect -798 712 -774 746
rect -740 712 -716 746
rect -798 674 -716 712
rect -798 640 -774 674
rect -740 640 -716 674
rect -798 602 -716 640
rect -798 568 -774 602
rect -740 568 -716 602
rect -798 530 -716 568
rect -798 496 -774 530
rect -740 496 -716 530
rect -798 458 -716 496
rect -798 424 -774 458
rect -740 424 -716 458
rect -798 386 -716 424
rect -798 352 -774 386
rect -740 352 -716 386
rect -798 314 -716 352
rect -798 280 -774 314
rect -740 280 -716 314
rect -798 242 -716 280
rect -798 208 -774 242
rect -740 208 -716 242
rect -798 170 -716 208
rect -798 136 -774 170
rect -740 136 -716 170
rect -798 98 -716 136
rect -798 64 -774 98
rect -740 64 -716 98
rect -798 26 -716 64
rect -798 -8 -774 26
rect -740 -8 -716 26
rect -798 -46 -716 -8
rect -798 -80 -774 -46
rect -740 -80 -716 -46
rect -798 -118 -716 -80
rect -798 -152 -774 -118
rect -740 -152 -716 -118
rect -798 -190 -716 -152
rect -659 6146 -457 6165
rect -659 6127 -647 6146
rect -469 6127 -457 6146
rect -659 -133 -648 6127
rect -468 -133 -457 6127
rect -659 -152 -647 -133
rect -469 -152 -457 -133
rect -659 -164 -457 -152
rect -134 6146 284 6165
rect -134 -152 -122 6146
rect 272 -152 284 6146
rect -134 -164 284 -152
rect 607 6146 809 6165
rect 607 6127 619 6146
rect 797 6127 809 6146
rect 607 -133 618 6127
rect 798 -133 809 6127
rect 607 -152 619 -133
rect 797 -152 809 -133
rect 607 -164 809 -152
rect 866 6146 948 6184
rect 866 6112 890 6146
rect 924 6112 948 6146
rect 866 6074 948 6112
rect 866 6040 890 6074
rect 924 6040 948 6074
rect 866 6002 948 6040
rect 866 5968 890 6002
rect 924 5968 948 6002
rect 866 5930 948 5968
rect 866 5896 890 5930
rect 924 5896 948 5930
rect 866 5858 948 5896
rect 866 5824 890 5858
rect 924 5824 948 5858
rect 866 5786 948 5824
rect 866 5752 890 5786
rect 924 5752 948 5786
rect 866 5714 948 5752
rect 866 5680 890 5714
rect 924 5680 948 5714
rect 866 5642 948 5680
rect 866 5608 890 5642
rect 924 5608 948 5642
rect 866 5570 948 5608
rect 866 5536 890 5570
rect 924 5536 948 5570
rect 866 5498 948 5536
rect 866 5464 890 5498
rect 924 5464 948 5498
rect 866 5426 948 5464
rect 866 5392 890 5426
rect 924 5392 948 5426
rect 866 5354 948 5392
rect 866 5320 890 5354
rect 924 5320 948 5354
rect 866 5282 948 5320
rect 866 5248 890 5282
rect 924 5248 948 5282
rect 866 5210 948 5248
rect 866 5176 890 5210
rect 924 5176 948 5210
rect 866 5138 948 5176
rect 866 5104 890 5138
rect 924 5104 948 5138
rect 866 5066 948 5104
rect 866 5032 890 5066
rect 924 5032 948 5066
rect 866 4994 948 5032
rect 866 4960 890 4994
rect 924 4960 948 4994
rect 866 4922 948 4960
rect 866 4888 890 4922
rect 924 4888 948 4922
rect 866 4850 948 4888
rect 866 4816 890 4850
rect 924 4816 948 4850
rect 866 4778 948 4816
rect 866 4744 890 4778
rect 924 4744 948 4778
rect 866 4706 948 4744
rect 866 4672 890 4706
rect 924 4672 948 4706
rect 866 4634 948 4672
rect 866 4600 890 4634
rect 924 4600 948 4634
rect 866 4562 948 4600
rect 866 4528 890 4562
rect 924 4528 948 4562
rect 866 4490 948 4528
rect 866 4456 890 4490
rect 924 4456 948 4490
rect 866 4418 948 4456
rect 866 4384 890 4418
rect 924 4384 948 4418
rect 866 4346 948 4384
rect 866 4312 890 4346
rect 924 4312 948 4346
rect 866 4274 948 4312
rect 866 4240 890 4274
rect 924 4240 948 4274
rect 866 4202 948 4240
rect 866 4168 890 4202
rect 924 4168 948 4202
rect 866 4130 948 4168
rect 866 4096 890 4130
rect 924 4096 948 4130
rect 866 4058 948 4096
rect 866 4024 890 4058
rect 924 4024 948 4058
rect 866 3986 948 4024
rect 866 3952 890 3986
rect 924 3952 948 3986
rect 866 3914 948 3952
rect 866 3880 890 3914
rect 924 3880 948 3914
rect 866 3842 948 3880
rect 866 3808 890 3842
rect 924 3808 948 3842
rect 866 3770 948 3808
rect 866 3736 890 3770
rect 924 3736 948 3770
rect 866 3698 948 3736
rect 866 3664 890 3698
rect 924 3664 948 3698
rect 866 3626 948 3664
rect 866 3592 890 3626
rect 924 3592 948 3626
rect 866 3554 948 3592
rect 866 3520 890 3554
rect 924 3520 948 3554
rect 866 3482 948 3520
rect 866 3448 890 3482
rect 924 3448 948 3482
rect 866 3410 948 3448
rect 866 3376 890 3410
rect 924 3376 948 3410
rect 866 3338 948 3376
rect 866 3304 890 3338
rect 924 3304 948 3338
rect 866 3266 948 3304
rect 866 3232 890 3266
rect 924 3232 948 3266
rect 866 3194 948 3232
rect 866 3160 890 3194
rect 924 3160 948 3194
rect 866 3122 948 3160
rect 866 3088 890 3122
rect 924 3088 948 3122
rect 866 3050 948 3088
rect 866 3016 890 3050
rect 924 3016 948 3050
rect 866 2978 948 3016
rect 866 2944 890 2978
rect 924 2944 948 2978
rect 866 2906 948 2944
rect 866 2872 890 2906
rect 924 2872 948 2906
rect 866 2834 948 2872
rect 866 2800 890 2834
rect 924 2800 948 2834
rect 866 2762 948 2800
rect 866 2728 890 2762
rect 924 2728 948 2762
rect 866 2690 948 2728
rect 866 2656 890 2690
rect 924 2656 948 2690
rect 866 2618 948 2656
rect 866 2584 890 2618
rect 924 2584 948 2618
rect 866 2546 948 2584
rect 866 2512 890 2546
rect 924 2512 948 2546
rect 866 2474 948 2512
rect 866 2440 890 2474
rect 924 2440 948 2474
rect 866 2402 948 2440
rect 866 2368 890 2402
rect 924 2368 948 2402
rect 866 2330 948 2368
rect 866 2296 890 2330
rect 924 2296 948 2330
rect 866 2258 948 2296
rect 866 2224 890 2258
rect 924 2224 948 2258
rect 866 2186 948 2224
rect 866 2152 890 2186
rect 924 2152 948 2186
rect 866 2114 948 2152
rect 866 2080 890 2114
rect 924 2080 948 2114
rect 866 2042 948 2080
rect 866 2008 890 2042
rect 924 2008 948 2042
rect 866 1970 948 2008
rect 866 1936 890 1970
rect 924 1936 948 1970
rect 866 1898 948 1936
rect 866 1864 890 1898
rect 924 1864 948 1898
rect 866 1826 948 1864
rect 866 1792 890 1826
rect 924 1792 948 1826
rect 866 1754 948 1792
rect 866 1720 890 1754
rect 924 1720 948 1754
rect 866 1682 948 1720
rect 866 1648 890 1682
rect 924 1648 948 1682
rect 866 1610 948 1648
rect 866 1576 890 1610
rect 924 1576 948 1610
rect 866 1538 948 1576
rect 866 1504 890 1538
rect 924 1504 948 1538
rect 866 1466 948 1504
rect 866 1432 890 1466
rect 924 1432 948 1466
rect 866 1394 948 1432
rect 866 1360 890 1394
rect 924 1360 948 1394
rect 866 1322 948 1360
rect 866 1288 890 1322
rect 924 1288 948 1322
rect 866 1250 948 1288
rect 866 1216 890 1250
rect 924 1216 948 1250
rect 866 1178 948 1216
rect 866 1144 890 1178
rect 924 1144 948 1178
rect 866 1106 948 1144
rect 866 1072 890 1106
rect 924 1072 948 1106
rect 866 1034 948 1072
rect 866 1000 890 1034
rect 924 1000 948 1034
rect 866 962 948 1000
rect 866 928 890 962
rect 924 928 948 962
rect 866 890 948 928
rect 866 856 890 890
rect 924 856 948 890
rect 866 818 948 856
rect 866 784 890 818
rect 924 784 948 818
rect 866 746 948 784
rect 866 712 890 746
rect 924 712 948 746
rect 866 674 948 712
rect 866 640 890 674
rect 924 640 948 674
rect 866 602 948 640
rect 866 568 890 602
rect 924 568 948 602
rect 866 530 948 568
rect 866 496 890 530
rect 924 496 948 530
rect 866 458 948 496
rect 866 424 890 458
rect 924 424 948 458
rect 866 386 948 424
rect 866 352 890 386
rect 924 352 948 386
rect 866 314 948 352
rect 866 280 890 314
rect 924 280 948 314
rect 866 242 948 280
rect 866 208 890 242
rect 924 208 948 242
rect 866 170 948 208
rect 866 136 890 170
rect 924 136 948 170
rect 866 98 948 136
rect 866 64 890 98
rect 924 64 948 98
rect 866 26 948 64
rect 866 -8 890 26
rect 924 -8 948 26
rect 866 -46 948 -8
rect 866 -80 890 -46
rect 924 -80 948 -46
rect 866 -118 948 -80
rect 866 -152 890 -118
rect 924 -152 948 -118
rect -798 -224 -774 -190
rect -740 -224 -716 -190
rect -798 -262 -716 -224
rect -798 -296 -774 -262
rect -740 -296 -716 -262
rect -798 -334 -716 -296
rect -798 -368 -774 -334
rect -740 -368 -716 -334
rect -798 -406 -716 -368
rect -798 -440 -774 -406
rect -740 -440 -716 -406
rect -798 -478 -716 -440
rect 866 -190 948 -152
rect 866 -224 890 -190
rect 924 -224 948 -190
rect 866 -262 948 -224
rect 866 -296 890 -262
rect 924 -296 948 -262
rect 866 -334 948 -296
rect 866 -368 890 -334
rect 924 -368 948 -334
rect 866 -406 948 -368
rect 866 -440 890 -406
rect 924 -440 948 -406
rect -798 -512 -774 -478
rect -740 -512 -716 -478
rect -798 -550 -716 -512
rect -798 -584 -774 -550
rect -740 -584 -716 -550
rect -798 -622 -716 -584
rect -798 -656 -774 -622
rect -740 -656 -716 -622
rect -798 -757 -716 -656
rect -146 -450 290 -443
rect -146 -502 -139 -450
rect -87 -502 -65 -450
rect -13 -502 9 -450
rect 61 -502 83 -450
rect 135 -502 157 -450
rect 209 -502 231 -450
rect 283 -502 290 -450
rect -146 -524 290 -502
rect -146 -576 -139 -524
rect -87 -576 -65 -524
rect -13 -576 9 -524
rect 61 -576 83 -524
rect 135 -576 157 -524
rect 209 -576 231 -524
rect 283 -576 290 -524
rect -146 -598 290 -576
rect -146 -650 -139 -598
rect -87 -650 -65 -598
rect -13 -650 9 -598
rect 61 -650 83 -598
rect 135 -650 157 -598
rect 209 -650 231 -598
rect 283 -650 290 -598
rect -146 -657 290 -650
rect 866 -478 948 -440
rect 866 -512 890 -478
rect 924 -512 948 -478
rect 866 -550 948 -512
rect 866 -584 890 -550
rect 924 -584 948 -550
rect 866 -622 948 -584
rect 866 -656 890 -622
rect 924 -656 948 -622
rect 866 -757 948 -656
rect -798 -820 948 -757
rect -798 -998 -554 -820
rect 704 -998 948 -820
rect -798 -1022 948 -998
rect 1648 7013 1730 7051
rect 1648 6979 1672 7013
rect 1706 6979 1730 7013
rect 1648 6941 1730 6979
rect 1648 6907 1672 6941
rect 1706 6907 1730 6941
rect 1648 6869 1730 6907
rect 1648 6835 1672 6869
rect 1706 6835 1730 6869
rect 1648 6797 1730 6835
rect 1648 6763 1672 6797
rect 1706 6763 1730 6797
rect 1648 6725 1730 6763
rect 1648 6691 1672 6725
rect 1706 6691 1730 6725
rect 1648 6653 1730 6691
rect 1648 6619 1672 6653
rect 1706 6619 1730 6653
rect 1648 6581 1730 6619
rect 1648 6547 1672 6581
rect 1706 6547 1730 6581
rect 1648 6509 1730 6547
rect 1648 6475 1672 6509
rect 1706 6475 1730 6509
rect 1648 6437 1730 6475
rect 1648 6403 1672 6437
rect 1706 6403 1730 6437
rect 1648 6365 1730 6403
rect 1648 6331 1672 6365
rect 1706 6331 1730 6365
rect 1648 6293 1730 6331
rect 1648 6259 1672 6293
rect 1706 6259 1730 6293
rect 1648 6221 1730 6259
rect 1648 6187 1672 6221
rect 1706 6187 1730 6221
rect 1648 6149 1730 6187
rect 1648 6115 1672 6149
rect 1706 6115 1730 6149
rect 1648 6077 1730 6115
rect 1648 6043 1672 6077
rect 1706 6043 1730 6077
rect 1648 6005 1730 6043
rect 1648 5971 1672 6005
rect 1706 5971 1730 6005
rect 1648 5933 1730 5971
rect 1648 5899 1672 5933
rect 1706 5899 1730 5933
rect 1648 5861 1730 5899
rect 1648 5827 1672 5861
rect 1706 5827 1730 5861
rect 1648 5789 1730 5827
rect 1648 5755 1672 5789
rect 1706 5755 1730 5789
rect 1648 5717 1730 5755
rect 1648 5683 1672 5717
rect 1706 5683 1730 5717
rect 1648 5645 1730 5683
rect 1648 5611 1672 5645
rect 1706 5611 1730 5645
rect 1648 5573 1730 5611
rect 1648 5539 1672 5573
rect 1706 5539 1730 5573
rect 1648 5501 1730 5539
rect 1648 5467 1672 5501
rect 1706 5467 1730 5501
rect 1648 5429 1730 5467
rect 1648 5395 1672 5429
rect 1706 5395 1730 5429
rect 1648 5357 1730 5395
rect 1648 5323 1672 5357
rect 1706 5323 1730 5357
rect 1648 5285 1730 5323
rect 1648 5251 1672 5285
rect 1706 5251 1730 5285
rect 1648 5213 1730 5251
rect 1648 5179 1672 5213
rect 1706 5179 1730 5213
rect 1648 5141 1730 5179
rect 1648 5107 1672 5141
rect 1706 5107 1730 5141
rect 1648 5069 1730 5107
rect 1648 5035 1672 5069
rect 1706 5035 1730 5069
rect 1648 4997 1730 5035
rect 1648 4963 1672 4997
rect 1706 4963 1730 4997
rect 1648 4925 1730 4963
rect 1648 4891 1672 4925
rect 1706 4891 1730 4925
rect 1648 4853 1730 4891
rect 1648 4819 1672 4853
rect 1706 4819 1730 4853
rect 1648 4781 1730 4819
rect 1648 4747 1672 4781
rect 1706 4747 1730 4781
rect 1648 4709 1730 4747
rect 1648 4675 1672 4709
rect 1706 4675 1730 4709
rect 1648 4637 1730 4675
rect 1648 4603 1672 4637
rect 1706 4603 1730 4637
rect 1648 4565 1730 4603
rect 1648 4531 1672 4565
rect 1706 4531 1730 4565
rect 1648 4493 1730 4531
rect 1648 4459 1672 4493
rect 1706 4459 1730 4493
rect 1648 4421 1730 4459
rect 1648 4387 1672 4421
rect 1706 4387 1730 4421
rect 1648 4349 1730 4387
rect 1648 4315 1672 4349
rect 1706 4315 1730 4349
rect 1648 4277 1730 4315
rect 1648 4243 1672 4277
rect 1706 4243 1730 4277
rect 1648 4205 1730 4243
rect 1648 4171 1672 4205
rect 1706 4171 1730 4205
rect 1648 4133 1730 4171
rect 1648 4099 1672 4133
rect 1706 4099 1730 4133
rect 1648 4061 1730 4099
rect 1648 4027 1672 4061
rect 1706 4027 1730 4061
rect 1648 3989 1730 4027
rect 1648 3955 1672 3989
rect 1706 3955 1730 3989
rect 1648 3917 1730 3955
rect 1648 3883 1672 3917
rect 1706 3883 1730 3917
rect 1648 3845 1730 3883
rect 1648 3811 1672 3845
rect 1706 3811 1730 3845
rect 1648 3773 1730 3811
rect 1648 3739 1672 3773
rect 1706 3739 1730 3773
rect 1648 3701 1730 3739
rect 1648 3667 1672 3701
rect 1706 3667 1730 3701
rect 1648 3629 1730 3667
rect 1648 3595 1672 3629
rect 1706 3595 1730 3629
rect 1648 3557 1730 3595
rect 1648 3523 1672 3557
rect 1706 3523 1730 3557
rect 1648 3485 1730 3523
rect 1648 3451 1672 3485
rect 1706 3451 1730 3485
rect 1648 3413 1730 3451
rect 1648 3379 1672 3413
rect 1706 3379 1730 3413
rect 1648 3341 1730 3379
rect 1648 3307 1672 3341
rect 1706 3307 1730 3341
rect 1648 3269 1730 3307
rect 1648 3235 1672 3269
rect 1706 3235 1730 3269
rect 1648 3197 1730 3235
rect 1648 3163 1672 3197
rect 1706 3163 1730 3197
rect 1648 3125 1730 3163
rect 1648 3091 1672 3125
rect 1706 3091 1730 3125
rect 1648 3053 1730 3091
rect 1648 3019 1672 3053
rect 1706 3019 1730 3053
rect 1648 2981 1730 3019
rect 1648 2947 1672 2981
rect 1706 2947 1730 2981
rect 1648 2909 1730 2947
rect 1648 2875 1672 2909
rect 1706 2875 1730 2909
rect 1648 2837 1730 2875
rect 1648 2803 1672 2837
rect 1706 2803 1730 2837
rect 1648 2765 1730 2803
rect 1648 2731 1672 2765
rect 1706 2731 1730 2765
rect 1648 2693 1730 2731
rect 1648 2659 1672 2693
rect 1706 2659 1730 2693
rect 1648 2621 1730 2659
rect 1648 2587 1672 2621
rect 1706 2587 1730 2621
rect 1648 2549 1730 2587
rect 1648 2515 1672 2549
rect 1706 2515 1730 2549
rect 1648 2477 1730 2515
rect 1648 2443 1672 2477
rect 1706 2443 1730 2477
rect 1648 2405 1730 2443
rect 1648 2371 1672 2405
rect 1706 2371 1730 2405
rect 1648 2333 1730 2371
rect 1648 2299 1672 2333
rect 1706 2299 1730 2333
rect 1648 2261 1730 2299
rect 1648 2227 1672 2261
rect 1706 2227 1730 2261
rect 1648 2189 1730 2227
rect 1648 2155 1672 2189
rect 1706 2155 1730 2189
rect 1648 2117 1730 2155
rect 1648 2083 1672 2117
rect 1706 2083 1730 2117
rect 1648 2045 1730 2083
rect 1648 2011 1672 2045
rect 1706 2011 1730 2045
rect 1648 1973 1730 2011
rect 1648 1939 1672 1973
rect 1706 1939 1730 1973
rect 1648 1901 1730 1939
rect 1648 1867 1672 1901
rect 1706 1867 1730 1901
rect 1648 1829 1730 1867
rect 1648 1795 1672 1829
rect 1706 1795 1730 1829
rect 1648 1757 1730 1795
rect 1648 1723 1672 1757
rect 1706 1723 1730 1757
rect 1648 1685 1730 1723
rect 1648 1651 1672 1685
rect 1706 1651 1730 1685
rect 1648 1613 1730 1651
rect 1648 1579 1672 1613
rect 1706 1579 1730 1613
rect 1648 1541 1730 1579
rect 1648 1507 1672 1541
rect 1706 1507 1730 1541
rect 1648 1469 1730 1507
rect 1648 1435 1672 1469
rect 1706 1435 1730 1469
rect 1648 1397 1730 1435
rect 1648 1363 1672 1397
rect 1706 1363 1730 1397
rect 1648 1325 1730 1363
rect 1648 1291 1672 1325
rect 1706 1291 1730 1325
rect 1648 1253 1730 1291
rect 1648 1219 1672 1253
rect 1706 1219 1730 1253
rect 1648 1181 1730 1219
rect 1648 1147 1672 1181
rect 1706 1147 1730 1181
rect 1648 1109 1730 1147
rect 1648 1075 1672 1109
rect 1706 1075 1730 1109
rect 1648 1037 1730 1075
rect 1648 1003 1672 1037
rect 1706 1003 1730 1037
rect 1648 965 1730 1003
rect 1648 931 1672 965
rect 1706 931 1730 965
rect 1648 893 1730 931
rect 1648 859 1672 893
rect 1706 859 1730 893
rect 1648 821 1730 859
rect 1648 787 1672 821
rect 1706 787 1730 821
rect 1648 749 1730 787
rect 1648 715 1672 749
rect 1706 715 1730 749
rect 1648 677 1730 715
rect 1648 643 1672 677
rect 1706 643 1730 677
rect 1648 605 1730 643
rect 1648 571 1672 605
rect 1706 571 1730 605
rect 1648 533 1730 571
rect 1648 499 1672 533
rect 1706 499 1730 533
rect 1648 461 1730 499
rect 1648 427 1672 461
rect 1706 427 1730 461
rect 1648 389 1730 427
rect 1648 355 1672 389
rect 1706 355 1730 389
rect 1648 317 1730 355
rect 1648 283 1672 317
rect 1706 283 1730 317
rect 1648 245 1730 283
rect 1648 211 1672 245
rect 1706 211 1730 245
rect 1648 173 1730 211
rect 1648 139 1672 173
rect 1706 139 1730 173
rect 1648 101 1730 139
rect 1648 67 1672 101
rect 1706 67 1730 101
rect 1648 29 1730 67
rect 1648 -5 1672 29
rect 1706 -5 1730 29
rect 1648 -43 1730 -5
rect 1648 -77 1672 -43
rect 1706 -77 1730 -43
rect 1648 -115 1730 -77
rect 1648 -149 1672 -115
rect 1706 -149 1730 -115
rect 1648 -187 1730 -149
rect 1648 -221 1672 -187
rect 1706 -221 1730 -187
rect 1648 -259 1730 -221
rect 1648 -293 1672 -259
rect 1706 -293 1730 -259
rect 1648 -331 1730 -293
rect 1648 -365 1672 -331
rect 1706 -365 1730 -331
rect 1648 -403 1730 -365
rect 1648 -437 1672 -403
rect 1706 -437 1730 -403
rect 1648 -475 1730 -437
rect 1648 -509 1672 -475
rect 1706 -509 1730 -475
rect 1648 -547 1730 -509
rect 1648 -581 1672 -547
rect 1706 -581 1730 -547
rect 1648 -619 1730 -581
rect 1648 -653 1672 -619
rect 1706 -653 1730 -619
rect 1648 -691 1730 -653
rect 1648 -725 1672 -691
rect 1706 -725 1730 -691
rect 1648 -763 1730 -725
rect 1648 -797 1672 -763
rect 1706 -797 1730 -763
rect 1648 -835 1730 -797
rect 1648 -869 1672 -835
rect 1706 -869 1730 -835
rect 1648 -907 1730 -869
rect 1648 -941 1672 -907
rect 1706 -941 1730 -907
rect 1648 -979 1730 -941
rect 1648 -1013 1672 -979
rect 1706 -1013 1730 -979
rect -1580 -1085 -1556 -1051
rect -1522 -1085 -1498 -1051
rect -1580 -1123 -1498 -1085
rect -1580 -1157 -1556 -1123
rect -1522 -1157 -1498 -1123
rect -1580 -1195 -1498 -1157
rect -1580 -1229 -1556 -1195
rect -1522 -1229 -1498 -1195
rect -1580 -1267 -1498 -1229
rect -1580 -1301 -1556 -1267
rect -1522 -1301 -1498 -1267
rect -1580 -1339 -1498 -1301
rect -1580 -1373 -1556 -1339
rect -1522 -1373 -1498 -1339
rect -1580 -1411 -1498 -1373
rect -1580 -1445 -1556 -1411
rect -1522 -1445 -1498 -1411
rect -1580 -1483 -1498 -1445
rect -1580 -1517 -1556 -1483
rect -1522 -1517 -1498 -1483
rect -1580 -1555 -1498 -1517
rect -1580 -1589 -1556 -1555
rect -1522 -1589 -1498 -1555
rect -1580 -1627 -1498 -1589
rect -1580 -1661 -1556 -1627
rect -1522 -1661 -1498 -1627
rect -1580 -1722 -1498 -1661
rect 1648 -1051 1730 -1013
rect 1648 -1085 1672 -1051
rect 1706 -1085 1730 -1051
rect 1648 -1123 1730 -1085
rect 1648 -1157 1672 -1123
rect 1706 -1157 1730 -1123
rect 1648 -1195 1730 -1157
rect 1648 -1229 1672 -1195
rect 1706 -1229 1730 -1195
rect 1648 -1267 1730 -1229
rect 1648 -1301 1672 -1267
rect 1706 -1301 1730 -1267
rect 1648 -1339 1730 -1301
rect 1648 -1373 1672 -1339
rect 1706 -1373 1730 -1339
rect 1648 -1411 1730 -1373
rect 1648 -1445 1672 -1411
rect 1706 -1445 1730 -1411
rect 1648 -1483 1730 -1445
rect 1648 -1517 1672 -1483
rect 1706 -1517 1730 -1483
rect 1648 -1555 1730 -1517
rect 1648 -1589 1672 -1555
rect 1706 -1589 1730 -1555
rect 1648 -1627 1730 -1589
rect 1648 -1661 1672 -1627
rect 1706 -1661 1730 -1627
rect 1648 -1722 1730 -1661
rect -1580 -1746 1730 -1722
rect -1580 -1780 -1454 -1746
rect -1420 -1780 -1382 -1746
rect -1348 -1780 -1310 -1746
rect -1276 -1780 -1238 -1746
rect -1204 -1780 -1166 -1746
rect -1132 -1780 -1094 -1746
rect -1060 -1780 -1022 -1746
rect -988 -1780 -950 -1746
rect -916 -1780 -878 -1746
rect -844 -1780 -806 -1746
rect -772 -1780 -734 -1746
rect -700 -1780 -662 -1746
rect -628 -1780 -590 -1746
rect -556 -1780 -518 -1746
rect -484 -1780 -446 -1746
rect -412 -1780 -374 -1746
rect -340 -1780 -302 -1746
rect -268 -1780 -230 -1746
rect -196 -1780 -158 -1746
rect -124 -1780 -86 -1746
rect -52 -1780 -14 -1746
rect 20 -1780 58 -1746
rect 92 -1780 130 -1746
rect 164 -1780 202 -1746
rect 236 -1780 274 -1746
rect 308 -1780 346 -1746
rect 380 -1780 418 -1746
rect 452 -1780 490 -1746
rect 524 -1780 562 -1746
rect 596 -1780 634 -1746
rect 668 -1780 706 -1746
rect 740 -1780 778 -1746
rect 812 -1780 850 -1746
rect 884 -1780 922 -1746
rect 956 -1780 994 -1746
rect 1028 -1780 1066 -1746
rect 1100 -1780 1138 -1746
rect 1172 -1780 1210 -1746
rect 1244 -1780 1282 -1746
rect 1316 -1780 1354 -1746
rect 1388 -1780 1426 -1746
rect 1460 -1780 1498 -1746
rect 1532 -1780 1570 -1746
rect 1604 -1780 1730 -1746
rect -1580 -1804 1730 -1780
<< via1 >>
rect -648 -133 -647 6127
rect -647 -133 -469 6127
rect -469 -133 -468 6127
rect -111 -133 261 6127
rect 618 -133 619 6127
rect 619 -133 797 6127
rect 797 -133 798 6127
rect -139 -459 -87 -450
rect -139 -493 -130 -459
rect -130 -493 -96 -459
rect -96 -493 -87 -459
rect -139 -502 -87 -493
rect -65 -459 -13 -450
rect -65 -493 -56 -459
rect -56 -493 -22 -459
rect -22 -493 -13 -459
rect -65 -502 -13 -493
rect 9 -459 61 -450
rect 9 -493 18 -459
rect 18 -493 52 -459
rect 52 -493 61 -459
rect 9 -502 61 -493
rect 83 -459 135 -450
rect 83 -493 92 -459
rect 92 -493 126 -459
rect 126 -493 135 -459
rect 83 -502 135 -493
rect 157 -459 209 -450
rect 157 -493 166 -459
rect 166 -493 200 -459
rect 200 -493 209 -459
rect 157 -502 209 -493
rect 231 -459 283 -450
rect 231 -493 240 -459
rect 240 -493 274 -459
rect 274 -493 283 -459
rect 231 -502 283 -493
rect -139 -533 -87 -524
rect -139 -567 -130 -533
rect -130 -567 -96 -533
rect -96 -567 -87 -533
rect -139 -576 -87 -567
rect -65 -533 -13 -524
rect -65 -567 -56 -533
rect -56 -567 -22 -533
rect -22 -567 -13 -533
rect -65 -576 -13 -567
rect 9 -533 61 -524
rect 9 -567 18 -533
rect 18 -567 52 -533
rect 52 -567 61 -533
rect 9 -576 61 -567
rect 83 -533 135 -524
rect 83 -567 92 -533
rect 92 -567 126 -533
rect 126 -567 135 -533
rect 83 -576 135 -567
rect 157 -533 209 -524
rect 157 -567 166 -533
rect 166 -567 200 -533
rect 200 -567 209 -533
rect 157 -576 209 -567
rect 231 -533 283 -524
rect 231 -567 240 -533
rect 240 -567 274 -533
rect 274 -567 283 -533
rect 231 -576 283 -567
rect -139 -607 -87 -598
rect -139 -641 -130 -607
rect -130 -641 -96 -607
rect -96 -641 -87 -607
rect -139 -650 -87 -641
rect -65 -607 -13 -598
rect -65 -641 -56 -607
rect -56 -641 -22 -607
rect -22 -641 -13 -607
rect -65 -650 -13 -641
rect 9 -607 61 -598
rect 9 -641 18 -607
rect 18 -641 52 -607
rect 52 -641 61 -607
rect 9 -650 61 -641
rect 83 -607 135 -598
rect 83 -641 92 -607
rect 92 -641 126 -607
rect 126 -641 135 -607
rect 83 -650 135 -641
rect 157 -607 209 -598
rect 157 -641 166 -607
rect 166 -641 200 -607
rect 200 -641 209 -607
rect 157 -650 209 -641
rect 231 -607 283 -598
rect 231 -641 240 -607
rect 240 -641 274 -607
rect 274 -641 283 -607
rect 231 -650 283 -641
<< metal2 >>
rect -659 6127 -457 6165
rect -659 -133 -648 6127
rect -468 -133 -457 6127
rect -659 -1122 -457 -133
rect -134 6127 284 7122
rect -134 -133 -111 6127
rect 261 -133 284 6127
rect -134 -164 284 -133
rect 607 6127 809 6165
rect 607 -133 618 6127
rect 798 -133 809 6127
rect -146 -450 290 -443
rect -146 -502 -139 -450
rect -87 -479 -65 -450
rect -13 -479 9 -450
rect 61 -479 83 -450
rect 135 -479 157 -450
rect 209 -479 231 -450
rect 283 -502 290 -450
rect -146 -524 -116 -502
rect 260 -524 290 -502
rect -146 -576 -139 -524
rect 283 -576 290 -524
rect -146 -598 -116 -576
rect 260 -598 290 -576
rect -146 -650 -139 -598
rect -87 -650 -65 -615
rect -13 -650 9 -615
rect 61 -650 83 -615
rect 135 -650 157 -615
rect 209 -650 231 -615
rect 283 -650 290 -598
rect -146 -657 290 -650
rect 607 -1122 809 -133
<< via2 >>
rect -116 -502 -87 -479
rect -87 -502 -65 -479
rect -65 -502 -13 -479
rect -13 -502 9 -479
rect 9 -502 61 -479
rect 61 -502 83 -479
rect 83 -502 135 -479
rect 135 -502 157 -479
rect 157 -502 209 -479
rect 209 -502 231 -479
rect 231 -502 260 -479
rect -116 -524 260 -502
rect -116 -576 -87 -524
rect -87 -576 -65 -524
rect -65 -576 -13 -524
rect -13 -576 9 -524
rect 9 -576 61 -524
rect 61 -576 83 -524
rect 83 -576 135 -524
rect 135 -576 157 -524
rect 157 -576 209 -524
rect 209 -576 231 -524
rect 231 -576 260 -524
rect -116 -598 260 -576
rect -116 -615 -87 -598
rect -87 -615 -65 -598
rect -65 -615 -13 -598
rect -13 -615 9 -598
rect 9 -615 61 -598
rect 61 -615 83 -598
rect 83 -615 135 -598
rect 135 -615 157 -598
rect 157 -615 209 -598
rect 209 -615 231 -598
rect 231 -615 260 -598
<< metal3 >>
rect -150 -479 290 -443
rect -150 -615 -116 -479
rect 260 -615 290 -479
rect -150 -657 290 -615
<< labels >>
flabel comment s 750 122 750 122 0 FreeSans 1600 0 0 0 S
flabel comment s -528 7380 -528 7380 0 FreeSans 1200 0 0 0 condiodeHvPsub
flabel comment s 62 122 62 122 0 FreeSans 1600 0 0 0 D
flabel comment s -589 122 -589 122 0 FreeSans 1600 0 0 0 S
<< properties >>
string GDS_END 10388286
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10116956
<< end >>
