magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 107 157 619 203
rect 1 21 735 157
rect 30 -17 64 21
<< scnmos >>
rect 81 47 111 131
rect 183 47 283 177
rect 443 47 543 177
rect 608 47 638 131
<< scpmoshvt >>
rect 81 297 111 497
rect 183 333 283 497
rect 443 333 543 497
rect 608 297 638 497
<< ndiff >>
rect 133 131 183 177
rect 27 104 81 131
rect 27 70 36 104
rect 70 70 81 104
rect 27 47 81 70
rect 111 104 183 131
rect 111 70 133 104
rect 167 70 183 104
rect 111 47 183 70
rect 283 104 335 177
rect 283 70 293 104
rect 327 70 335 104
rect 283 47 335 70
rect 390 104 443 177
rect 390 70 398 104
rect 432 70 443 104
rect 390 47 443 70
rect 543 131 593 177
rect 543 104 608 131
rect 543 70 554 104
rect 588 70 608 104
rect 543 47 608 70
rect 638 104 709 131
rect 638 70 652 104
rect 686 70 709 104
rect 638 47 709 70
<< pdiff >>
rect 27 478 81 497
rect 27 444 36 478
rect 70 444 81 478
rect 27 410 81 444
rect 27 376 36 410
rect 70 376 81 410
rect 27 297 81 376
rect 111 478 183 497
rect 111 444 136 478
rect 170 444 183 478
rect 111 410 183 444
rect 111 376 136 410
rect 170 376 183 410
rect 111 333 183 376
rect 283 478 336 497
rect 283 444 294 478
rect 328 444 336 478
rect 283 410 336 444
rect 283 376 294 410
rect 328 376 336 410
rect 283 333 336 376
rect 390 477 443 497
rect 390 443 398 477
rect 432 443 443 477
rect 390 409 443 443
rect 390 375 398 409
rect 432 375 443 409
rect 390 333 443 375
rect 543 478 608 497
rect 543 444 554 478
rect 588 444 608 478
rect 543 410 608 444
rect 543 376 554 410
rect 588 376 608 410
rect 543 333 608 376
rect 111 297 161 333
rect 558 297 608 333
rect 638 477 709 497
rect 638 443 652 477
rect 686 443 709 477
rect 638 409 709 443
rect 638 375 652 409
rect 686 375 709 409
rect 638 297 709 375
<< ndiffc >>
rect 36 70 70 104
rect 133 70 167 104
rect 293 70 327 104
rect 398 70 432 104
rect 554 70 588 104
rect 652 70 686 104
<< pdiffc >>
rect 36 444 70 478
rect 36 376 70 410
rect 136 444 170 478
rect 136 376 170 410
rect 294 444 328 478
rect 294 376 328 410
rect 398 443 432 477
rect 398 375 432 409
rect 554 444 588 478
rect 554 376 588 410
rect 652 443 686 477
rect 652 375 686 409
<< poly >>
rect 81 497 111 523
rect 183 497 283 523
rect 443 497 543 523
rect 608 497 638 523
rect 81 262 111 297
rect 41 249 111 262
rect 183 259 283 333
rect 443 259 543 333
rect 608 265 638 297
rect 41 215 57 249
rect 91 215 111 249
rect 41 203 111 215
rect 161 249 283 259
rect 161 215 177 249
rect 211 215 283 249
rect 161 205 283 215
rect 382 249 543 259
rect 382 215 398 249
rect 432 215 543 249
rect 382 205 543 215
rect 81 131 111 203
rect 183 177 283 205
rect 443 177 543 205
rect 588 249 642 265
rect 588 215 598 249
rect 632 215 642 249
rect 588 199 642 215
rect 608 131 638 199
rect 81 21 111 47
rect 183 21 283 47
rect 443 21 543 47
rect 608 21 638 47
<< polycont >>
rect 57 215 91 249
rect 177 215 211 249
rect 398 215 432 249
rect 598 215 632 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 478 86 493
rect 17 444 36 478
rect 70 444 86 478
rect 17 410 86 444
rect 17 376 36 410
rect 70 376 86 410
rect 17 326 86 376
rect 120 478 186 527
rect 120 444 136 478
rect 170 444 186 478
rect 120 410 186 444
rect 120 376 136 410
rect 170 376 186 410
rect 120 360 186 376
rect 276 478 346 493
rect 276 444 294 478
rect 328 444 346 478
rect 276 410 346 444
rect 276 376 294 410
rect 328 376 346 410
rect 17 292 211 326
rect 141 263 211 292
rect 276 264 346 376
rect 398 477 448 493
rect 432 443 448 477
rect 398 409 448 443
rect 432 375 448 409
rect 398 333 448 375
rect 538 478 604 527
rect 538 444 554 478
rect 588 444 604 478
rect 538 410 604 444
rect 538 376 554 410
rect 588 376 604 410
rect 538 367 604 376
rect 638 477 719 493
rect 638 443 652 477
rect 686 443 719 477
rect 638 409 719 443
rect 638 375 652 409
rect 686 375 719 409
rect 638 338 719 375
rect 398 299 516 333
rect 482 265 516 299
rect 17 249 107 258
rect 17 215 57 249
rect 91 215 107 249
rect 141 249 227 263
rect 141 215 177 249
rect 211 215 227 249
rect 141 205 227 215
rect 276 249 448 264
rect 276 215 398 249
rect 432 215 448 249
rect 276 214 448 215
rect 482 249 635 265
rect 482 215 598 249
rect 632 215 635 249
rect 141 181 211 205
rect 17 147 211 181
rect 17 104 83 147
rect 17 70 36 104
rect 70 70 83 104
rect 17 51 83 70
rect 117 104 183 113
rect 117 70 133 104
rect 167 70 183 104
rect 117 17 183 70
rect 276 104 346 214
rect 482 199 635 215
rect 482 180 516 199
rect 276 70 293 104
rect 327 70 346 104
rect 276 51 346 70
rect 398 146 516 180
rect 398 104 448 146
rect 669 128 719 338
rect 432 70 448 104
rect 398 51 448 70
rect 538 104 604 120
rect 538 70 554 104
rect 588 70 604 104
rect 538 17 604 70
rect 638 104 719 128
rect 638 70 652 104
rect 686 70 719 104
rect 638 51 719 70
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 676 425 710 459 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 676 357 710 391 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 676 289 710 323 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 676 221 710 255 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 676 153 710 187 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel locali s 676 85 710 119 0 FreeSans 400 0 0 0 X
port 6 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 clkdlybuf4s50_1
rlabel metal1 s 0 -48 736 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 736 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string GDS_END 3297142
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3290990
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 18.400 0.000 
<< end >>
