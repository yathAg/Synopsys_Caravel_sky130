magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect 0 0 776 1214
<< pmos >>
rect 204 102 254 1112
rect 310 102 360 1112
rect 416 102 466 1112
rect 522 102 572 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 254 1100 310 1112
rect 254 1066 265 1100
rect 299 1066 310 1100
rect 254 1032 310 1066
rect 254 998 265 1032
rect 299 998 310 1032
rect 254 964 310 998
rect 254 930 265 964
rect 299 930 310 964
rect 254 896 310 930
rect 254 862 265 896
rect 299 862 310 896
rect 254 828 310 862
rect 254 794 265 828
rect 299 794 310 828
rect 254 760 310 794
rect 254 726 265 760
rect 299 726 310 760
rect 254 692 310 726
rect 254 658 265 692
rect 299 658 310 692
rect 254 624 310 658
rect 254 590 265 624
rect 299 590 310 624
rect 254 556 310 590
rect 254 522 265 556
rect 299 522 310 556
rect 254 488 310 522
rect 254 454 265 488
rect 299 454 310 488
rect 254 420 310 454
rect 254 386 265 420
rect 299 386 310 420
rect 254 352 310 386
rect 254 318 265 352
rect 299 318 310 352
rect 254 284 310 318
rect 254 250 265 284
rect 299 250 310 284
rect 254 216 310 250
rect 254 182 265 216
rect 299 182 310 216
rect 254 148 310 182
rect 254 114 265 148
rect 299 114 310 148
rect 254 102 310 114
rect 360 1100 416 1112
rect 360 1066 371 1100
rect 405 1066 416 1100
rect 360 1032 416 1066
rect 360 998 371 1032
rect 405 998 416 1032
rect 360 964 416 998
rect 360 930 371 964
rect 405 930 416 964
rect 360 896 416 930
rect 360 862 371 896
rect 405 862 416 896
rect 360 828 416 862
rect 360 794 371 828
rect 405 794 416 828
rect 360 760 416 794
rect 360 726 371 760
rect 405 726 416 760
rect 360 692 416 726
rect 360 658 371 692
rect 405 658 416 692
rect 360 624 416 658
rect 360 590 371 624
rect 405 590 416 624
rect 360 556 416 590
rect 360 522 371 556
rect 405 522 416 556
rect 360 488 416 522
rect 360 454 371 488
rect 405 454 416 488
rect 360 420 416 454
rect 360 386 371 420
rect 405 386 416 420
rect 360 352 416 386
rect 360 318 371 352
rect 405 318 416 352
rect 360 284 416 318
rect 360 250 371 284
rect 405 250 416 284
rect 360 216 416 250
rect 360 182 371 216
rect 405 182 416 216
rect 360 148 416 182
rect 360 114 371 148
rect 405 114 416 148
rect 360 102 416 114
rect 466 1100 522 1112
rect 466 1066 477 1100
rect 511 1066 522 1100
rect 466 1032 522 1066
rect 466 998 477 1032
rect 511 998 522 1032
rect 466 964 522 998
rect 466 930 477 964
rect 511 930 522 964
rect 466 896 522 930
rect 466 862 477 896
rect 511 862 522 896
rect 466 828 522 862
rect 466 794 477 828
rect 511 794 522 828
rect 466 760 522 794
rect 466 726 477 760
rect 511 726 522 760
rect 466 692 522 726
rect 466 658 477 692
rect 511 658 522 692
rect 466 624 522 658
rect 466 590 477 624
rect 511 590 522 624
rect 466 556 522 590
rect 466 522 477 556
rect 511 522 522 556
rect 466 488 522 522
rect 466 454 477 488
rect 511 454 522 488
rect 466 420 522 454
rect 466 386 477 420
rect 511 386 522 420
rect 466 352 522 386
rect 466 318 477 352
rect 511 318 522 352
rect 466 284 522 318
rect 466 250 477 284
rect 511 250 522 284
rect 466 216 522 250
rect 466 182 477 216
rect 511 182 522 216
rect 466 148 522 182
rect 466 114 477 148
rect 511 114 522 148
rect 466 102 522 114
rect 572 1100 628 1112
rect 572 1066 583 1100
rect 617 1066 628 1100
rect 572 1032 628 1066
rect 572 998 583 1032
rect 617 998 628 1032
rect 572 964 628 998
rect 572 930 583 964
rect 617 930 628 964
rect 572 896 628 930
rect 572 862 583 896
rect 617 862 628 896
rect 572 828 628 862
rect 572 794 583 828
rect 617 794 628 828
rect 572 760 628 794
rect 572 726 583 760
rect 617 726 628 760
rect 572 692 628 726
rect 572 658 583 692
rect 617 658 628 692
rect 572 624 628 658
rect 572 590 583 624
rect 617 590 628 624
rect 572 556 628 590
rect 572 522 583 556
rect 617 522 628 556
rect 572 488 628 522
rect 572 454 583 488
rect 617 454 628 488
rect 572 420 628 454
rect 572 386 583 420
rect 617 386 628 420
rect 572 352 628 386
rect 572 318 583 352
rect 617 318 628 352
rect 572 284 628 318
rect 572 250 583 284
rect 617 250 628 284
rect 572 216 628 250
rect 572 182 583 216
rect 617 182 628 216
rect 572 148 628 182
rect 572 114 583 148
rect 617 114 628 148
rect 572 102 628 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 265 1066 299 1100
rect 265 998 299 1032
rect 265 930 299 964
rect 265 862 299 896
rect 265 794 299 828
rect 265 726 299 760
rect 265 658 299 692
rect 265 590 299 624
rect 265 522 299 556
rect 265 454 299 488
rect 265 386 299 420
rect 265 318 299 352
rect 265 250 299 284
rect 265 182 299 216
rect 265 114 299 148
rect 371 1066 405 1100
rect 371 998 405 1032
rect 371 930 405 964
rect 371 862 405 896
rect 371 794 405 828
rect 371 726 405 760
rect 371 658 405 692
rect 371 590 405 624
rect 371 522 405 556
rect 371 454 405 488
rect 371 386 405 420
rect 371 318 405 352
rect 371 250 405 284
rect 371 182 405 216
rect 371 114 405 148
rect 477 1066 511 1100
rect 477 998 511 1032
rect 477 930 511 964
rect 477 862 511 896
rect 477 794 511 828
rect 477 726 511 760
rect 477 658 511 692
rect 477 590 511 624
rect 477 522 511 556
rect 477 454 511 488
rect 477 386 511 420
rect 477 318 511 352
rect 477 250 511 284
rect 477 182 511 216
rect 477 114 511 148
rect 583 1066 617 1100
rect 583 998 617 1032
rect 583 930 617 964
rect 583 862 617 896
rect 583 794 617 828
rect 583 726 617 760
rect 583 658 617 692
rect 583 590 617 624
rect 583 522 617 556
rect 583 454 617 488
rect 583 386 617 420
rect 583 318 617 352
rect 583 250 617 284
rect 583 182 617 216
rect 583 114 617 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 682 1066 740 1112
rect 682 1032 694 1066
rect 728 1032 740 1066
rect 682 998 740 1032
rect 682 964 694 998
rect 728 964 740 998
rect 682 930 740 964
rect 682 896 694 930
rect 728 896 740 930
rect 682 862 740 896
rect 682 828 694 862
rect 728 828 740 862
rect 682 794 740 828
rect 682 760 694 794
rect 728 760 740 794
rect 682 726 740 760
rect 682 692 694 726
rect 728 692 740 726
rect 682 658 740 692
rect 682 624 694 658
rect 728 624 740 658
rect 682 590 740 624
rect 682 556 694 590
rect 728 556 740 590
rect 682 522 740 556
rect 682 488 694 522
rect 728 488 740 522
rect 682 454 740 488
rect 682 420 694 454
rect 728 420 740 454
rect 682 386 740 420
rect 682 352 694 386
rect 728 352 740 386
rect 682 318 740 352
rect 682 284 694 318
rect 728 284 740 318
rect 682 250 740 284
rect 682 216 694 250
rect 728 216 740 250
rect 682 182 740 216
rect 682 148 694 182
rect 728 148 740 182
rect 682 102 740 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 694 1032 728 1066
rect 694 964 728 998
rect 694 896 728 930
rect 694 828 728 862
rect 694 760 728 794
rect 694 692 728 726
rect 694 624 728 658
rect 694 556 728 590
rect 694 488 728 522
rect 694 420 728 454
rect 694 352 728 386
rect 694 284 728 318
rect 694 216 728 250
rect 694 148 728 182
<< poly >>
rect 185 1194 591 1214
rect 185 1160 201 1194
rect 235 1160 269 1194
rect 303 1160 337 1194
rect 371 1160 405 1194
rect 439 1160 473 1194
rect 507 1160 541 1194
rect 575 1160 591 1194
rect 185 1144 591 1160
rect 204 1112 254 1144
rect 310 1112 360 1144
rect 416 1112 466 1144
rect 522 1112 572 1144
rect 204 70 254 102
rect 310 70 360 102
rect 416 70 466 102
rect 522 70 572 102
rect 185 54 591 70
rect 185 20 201 54
rect 235 20 269 54
rect 303 20 337 54
rect 371 20 405 54
rect 439 20 473 54
rect 507 20 541 54
rect 575 20 591 54
rect 185 0 591 20
<< polycont >>
rect 201 1160 235 1194
rect 269 1160 303 1194
rect 337 1160 371 1194
rect 405 1160 439 1194
rect 473 1160 507 1194
rect 541 1160 575 1194
rect 201 20 235 54
rect 269 20 303 54
rect 337 20 371 54
rect 405 20 439 54
rect 473 20 507 54
rect 541 20 575 54
<< locali >>
rect 185 1160 192 1194
rect 235 1160 264 1194
rect 303 1160 336 1194
rect 371 1160 405 1194
rect 442 1160 473 1194
rect 514 1160 541 1194
rect 586 1160 591 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 265 1100 299 1116
rect 265 1032 299 1058
rect 265 964 299 986
rect 265 896 299 914
rect 265 828 299 842
rect 265 760 299 770
rect 265 692 299 698
rect 265 624 299 626
rect 265 588 299 590
rect 265 516 299 522
rect 265 444 299 454
rect 265 372 299 386
rect 265 300 299 318
rect 265 228 299 250
rect 265 156 299 182
rect 265 98 299 114
rect 371 1100 405 1116
rect 371 1032 405 1058
rect 371 964 405 986
rect 371 896 405 914
rect 371 828 405 842
rect 371 760 405 770
rect 371 692 405 698
rect 371 624 405 626
rect 371 588 405 590
rect 371 516 405 522
rect 371 444 405 454
rect 371 372 405 386
rect 371 300 405 318
rect 371 228 405 250
rect 371 156 405 182
rect 371 98 405 114
rect 477 1100 511 1116
rect 477 1032 511 1058
rect 477 964 511 986
rect 477 896 511 914
rect 477 828 511 842
rect 477 760 511 770
rect 477 692 511 698
rect 477 624 511 626
rect 477 588 511 590
rect 477 516 511 522
rect 477 444 511 454
rect 477 372 511 386
rect 477 300 511 318
rect 477 228 511 250
rect 477 156 511 182
rect 477 98 511 114
rect 583 1100 617 1116
rect 583 1032 617 1058
rect 583 964 617 986
rect 583 896 617 914
rect 583 828 617 842
rect 583 760 617 770
rect 583 692 617 698
rect 583 624 617 626
rect 583 588 617 590
rect 583 516 617 522
rect 583 444 617 454
rect 583 372 617 386
rect 583 300 617 318
rect 583 228 617 250
rect 583 156 617 182
rect 694 1020 728 1032
rect 694 948 728 964
rect 694 876 728 896
rect 694 804 728 828
rect 694 732 728 760
rect 694 660 728 692
rect 694 590 728 624
rect 694 522 728 554
rect 694 454 728 482
rect 694 386 728 410
rect 694 318 728 338
rect 694 250 728 266
rect 694 182 728 194
rect 583 98 617 114
rect 185 20 192 54
rect 235 20 264 54
rect 303 20 336 54
rect 371 20 405 54
rect 442 20 473 54
rect 514 20 541 54
rect 586 20 591 54
<< viali >>
rect 192 1160 201 1194
rect 201 1160 226 1194
rect 264 1160 269 1194
rect 269 1160 298 1194
rect 336 1160 337 1194
rect 337 1160 370 1194
rect 408 1160 439 1194
rect 439 1160 442 1194
rect 480 1160 507 1194
rect 507 1160 514 1194
rect 552 1160 575 1194
rect 575 1160 586 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 265 1066 299 1092
rect 265 1058 299 1066
rect 265 998 299 1020
rect 265 986 299 998
rect 265 930 299 948
rect 265 914 299 930
rect 265 862 299 876
rect 265 842 299 862
rect 265 794 299 804
rect 265 770 299 794
rect 265 726 299 732
rect 265 698 299 726
rect 265 658 299 660
rect 265 626 299 658
rect 265 556 299 588
rect 265 554 299 556
rect 265 488 299 516
rect 265 482 299 488
rect 265 420 299 444
rect 265 410 299 420
rect 265 352 299 372
rect 265 338 299 352
rect 265 284 299 300
rect 265 266 299 284
rect 265 216 299 228
rect 265 194 299 216
rect 265 148 299 156
rect 265 122 299 148
rect 371 1066 405 1092
rect 371 1058 405 1066
rect 371 998 405 1020
rect 371 986 405 998
rect 371 930 405 948
rect 371 914 405 930
rect 371 862 405 876
rect 371 842 405 862
rect 371 794 405 804
rect 371 770 405 794
rect 371 726 405 732
rect 371 698 405 726
rect 371 658 405 660
rect 371 626 405 658
rect 371 556 405 588
rect 371 554 405 556
rect 371 488 405 516
rect 371 482 405 488
rect 371 420 405 444
rect 371 410 405 420
rect 371 352 405 372
rect 371 338 405 352
rect 371 284 405 300
rect 371 266 405 284
rect 371 216 405 228
rect 371 194 405 216
rect 371 148 405 156
rect 371 122 405 148
rect 477 1066 511 1092
rect 477 1058 511 1066
rect 477 998 511 1020
rect 477 986 511 998
rect 477 930 511 948
rect 477 914 511 930
rect 477 862 511 876
rect 477 842 511 862
rect 477 794 511 804
rect 477 770 511 794
rect 477 726 511 732
rect 477 698 511 726
rect 477 658 511 660
rect 477 626 511 658
rect 477 556 511 588
rect 477 554 511 556
rect 477 488 511 516
rect 477 482 511 488
rect 477 420 511 444
rect 477 410 511 420
rect 477 352 511 372
rect 477 338 511 352
rect 477 284 511 300
rect 477 266 511 284
rect 477 216 511 228
rect 477 194 511 216
rect 477 148 511 156
rect 477 122 511 148
rect 583 1066 617 1092
rect 583 1058 617 1066
rect 583 998 617 1020
rect 583 986 617 998
rect 583 930 617 948
rect 583 914 617 930
rect 583 862 617 876
rect 583 842 617 862
rect 583 794 617 804
rect 583 770 617 794
rect 583 726 617 732
rect 583 698 617 726
rect 583 658 617 660
rect 583 626 617 658
rect 583 556 617 588
rect 583 554 617 556
rect 583 488 617 516
rect 583 482 617 488
rect 583 420 617 444
rect 583 410 617 420
rect 583 352 617 372
rect 583 338 617 352
rect 583 284 617 300
rect 583 266 617 284
rect 583 216 617 228
rect 583 194 617 216
rect 583 148 617 156
rect 583 122 617 148
rect 694 1066 728 1092
rect 694 1058 728 1066
rect 694 998 728 1020
rect 694 986 728 998
rect 694 930 728 948
rect 694 914 728 930
rect 694 862 728 876
rect 694 842 728 862
rect 694 794 728 804
rect 694 770 728 794
rect 694 726 728 732
rect 694 698 728 726
rect 694 658 728 660
rect 694 626 728 658
rect 694 556 728 588
rect 694 554 728 556
rect 694 488 728 516
rect 694 482 728 488
rect 694 420 728 444
rect 694 410 728 420
rect 694 352 728 372
rect 694 338 728 352
rect 694 284 728 300
rect 694 266 728 284
rect 694 216 728 228
rect 694 194 728 216
rect 694 148 728 156
rect 694 122 728 148
rect 192 20 201 54
rect 201 20 226 54
rect 264 20 269 54
rect 269 20 298 54
rect 336 20 337 54
rect 337 20 370 54
rect 408 20 439 54
rect 439 20 442 54
rect 480 20 507 54
rect 507 20 514 54
rect 552 20 575 54
rect 575 20 586 54
<< metal1 >>
rect 180 1194 598 1214
rect 180 1160 192 1194
rect 226 1160 264 1194
rect 298 1160 336 1194
rect 370 1160 408 1194
rect 442 1160 480 1194
rect 514 1160 552 1194
rect 586 1160 598 1194
rect 180 1148 598 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 256 1098 308 1104
rect 256 1034 308 1046
rect 256 970 308 982
rect 256 914 265 918
rect 299 914 308 918
rect 256 906 308 914
rect 256 842 265 854
rect 299 842 308 854
rect 256 778 265 790
rect 299 778 308 790
rect 256 714 265 726
rect 299 714 308 726
rect 256 660 308 662
rect 256 626 265 660
rect 299 626 308 660
rect 256 588 308 626
rect 256 554 265 588
rect 299 554 308 588
rect 256 516 308 554
rect 256 482 265 516
rect 299 482 308 516
rect 256 444 308 482
rect 256 410 265 444
rect 299 410 308 444
rect 256 372 308 410
rect 256 338 265 372
rect 299 338 308 372
rect 256 300 308 338
rect 256 266 265 300
rect 299 266 308 300
rect 256 228 308 266
rect 256 194 265 228
rect 299 194 308 228
rect 256 156 308 194
rect 256 122 265 156
rect 299 122 308 156
rect 256 110 308 122
rect 362 1092 414 1104
rect 362 1058 371 1092
rect 405 1058 414 1092
rect 362 1020 414 1058
rect 362 986 371 1020
rect 405 986 414 1020
rect 362 948 414 986
rect 362 914 371 948
rect 405 914 414 948
rect 362 876 414 914
rect 362 842 371 876
rect 405 842 414 876
rect 362 804 414 842
rect 362 770 371 804
rect 405 770 414 804
rect 362 732 414 770
rect 362 698 371 732
rect 405 698 414 732
rect 362 660 414 698
rect 362 626 371 660
rect 405 626 414 660
rect 362 588 414 626
rect 362 554 371 588
rect 405 554 414 588
rect 362 552 414 554
rect 362 488 371 500
rect 405 488 414 500
rect 362 424 371 436
rect 405 424 414 436
rect 362 360 371 372
rect 405 360 414 372
rect 362 300 414 308
rect 362 296 371 300
rect 405 296 414 300
rect 362 232 414 244
rect 362 168 414 180
rect 362 110 414 116
rect 468 1098 520 1104
rect 468 1034 520 1046
rect 468 970 520 982
rect 468 914 477 918
rect 511 914 520 918
rect 468 906 520 914
rect 468 842 477 854
rect 511 842 520 854
rect 468 778 477 790
rect 511 778 520 790
rect 468 714 477 726
rect 511 714 520 726
rect 468 660 520 662
rect 468 626 477 660
rect 511 626 520 660
rect 468 588 520 626
rect 468 554 477 588
rect 511 554 520 588
rect 468 516 520 554
rect 468 482 477 516
rect 511 482 520 516
rect 468 444 520 482
rect 468 410 477 444
rect 511 410 520 444
rect 468 372 520 410
rect 468 338 477 372
rect 511 338 520 372
rect 468 300 520 338
rect 468 266 477 300
rect 511 266 520 300
rect 468 228 520 266
rect 468 194 477 228
rect 511 194 520 228
rect 468 156 520 194
rect 468 122 477 156
rect 511 122 520 156
rect 468 110 520 122
rect 574 1092 626 1104
rect 574 1058 583 1092
rect 617 1058 626 1092
rect 574 1020 626 1058
rect 574 986 583 1020
rect 617 986 626 1020
rect 574 948 626 986
rect 574 914 583 948
rect 617 914 626 948
rect 574 876 626 914
rect 574 842 583 876
rect 617 842 626 876
rect 574 804 626 842
rect 574 770 583 804
rect 617 770 626 804
rect 574 732 626 770
rect 574 698 583 732
rect 617 698 626 732
rect 574 660 626 698
rect 574 626 583 660
rect 617 626 626 660
rect 574 588 626 626
rect 574 554 583 588
rect 617 554 626 588
rect 574 552 626 554
rect 574 488 583 500
rect 617 488 626 500
rect 574 424 583 436
rect 617 424 626 436
rect 574 360 583 372
rect 617 360 626 372
rect 574 300 626 308
rect 574 296 583 300
rect 617 296 626 300
rect 574 232 626 244
rect 574 168 626 180
rect 574 110 626 116
rect 682 1092 740 1104
rect 682 1058 694 1092
rect 728 1058 740 1092
rect 682 1020 740 1058
rect 682 986 694 1020
rect 728 986 740 1020
rect 682 948 740 986
rect 682 914 694 948
rect 728 914 740 948
rect 682 876 740 914
rect 682 842 694 876
rect 728 842 740 876
rect 682 804 740 842
rect 682 770 694 804
rect 728 770 740 804
rect 682 732 740 770
rect 682 698 694 732
rect 728 698 740 732
rect 682 660 740 698
rect 682 626 694 660
rect 728 626 740 660
rect 682 588 740 626
rect 682 554 694 588
rect 728 554 740 588
rect 682 516 740 554
rect 682 482 694 516
rect 728 482 740 516
rect 682 444 740 482
rect 682 410 694 444
rect 728 410 740 444
rect 682 372 740 410
rect 682 338 694 372
rect 728 338 740 372
rect 682 300 740 338
rect 682 266 694 300
rect 728 266 740 300
rect 682 228 740 266
rect 682 194 694 228
rect 728 194 740 228
rect 682 156 740 194
rect 682 122 694 156
rect 728 122 740 156
rect 682 110 740 122
rect 180 54 598 66
rect 180 20 192 54
rect 226 20 264 54
rect 298 20 336 54
rect 370 20 408 54
rect 442 20 480 54
rect 514 20 552 54
rect 586 20 598 54
rect 180 0 598 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 256 1092 308 1098
rect 256 1058 265 1092
rect 265 1058 299 1092
rect 299 1058 308 1092
rect 256 1046 308 1058
rect 256 1020 308 1034
rect 256 986 265 1020
rect 265 986 299 1020
rect 299 986 308 1020
rect 256 982 308 986
rect 256 948 308 970
rect 256 918 265 948
rect 265 918 299 948
rect 299 918 308 948
rect 256 876 308 906
rect 256 854 265 876
rect 265 854 299 876
rect 299 854 308 876
rect 256 804 308 842
rect 256 790 265 804
rect 265 790 299 804
rect 299 790 308 804
rect 256 770 265 778
rect 265 770 299 778
rect 299 770 308 778
rect 256 732 308 770
rect 256 726 265 732
rect 265 726 299 732
rect 299 726 308 732
rect 256 698 265 714
rect 265 698 299 714
rect 299 698 308 714
rect 256 662 308 698
rect 362 516 414 552
rect 362 500 371 516
rect 371 500 405 516
rect 405 500 414 516
rect 362 482 371 488
rect 371 482 405 488
rect 405 482 414 488
rect 362 444 414 482
rect 362 436 371 444
rect 371 436 405 444
rect 405 436 414 444
rect 362 410 371 424
rect 371 410 405 424
rect 405 410 414 424
rect 362 372 414 410
rect 362 338 371 360
rect 371 338 405 360
rect 405 338 414 360
rect 362 308 414 338
rect 362 266 371 296
rect 371 266 405 296
rect 405 266 414 296
rect 362 244 414 266
rect 362 228 414 232
rect 362 194 371 228
rect 371 194 405 228
rect 405 194 414 228
rect 362 180 414 194
rect 362 156 414 168
rect 362 122 371 156
rect 371 122 405 156
rect 405 122 414 156
rect 362 116 414 122
rect 468 1092 520 1098
rect 468 1058 477 1092
rect 477 1058 511 1092
rect 511 1058 520 1092
rect 468 1046 520 1058
rect 468 1020 520 1034
rect 468 986 477 1020
rect 477 986 511 1020
rect 511 986 520 1020
rect 468 982 520 986
rect 468 948 520 970
rect 468 918 477 948
rect 477 918 511 948
rect 511 918 520 948
rect 468 876 520 906
rect 468 854 477 876
rect 477 854 511 876
rect 511 854 520 876
rect 468 804 520 842
rect 468 790 477 804
rect 477 790 511 804
rect 511 790 520 804
rect 468 770 477 778
rect 477 770 511 778
rect 511 770 520 778
rect 468 732 520 770
rect 468 726 477 732
rect 477 726 511 732
rect 511 726 520 732
rect 468 698 477 714
rect 477 698 511 714
rect 511 698 520 714
rect 468 662 520 698
rect 574 516 626 552
rect 574 500 583 516
rect 583 500 617 516
rect 617 500 626 516
rect 574 482 583 488
rect 583 482 617 488
rect 617 482 626 488
rect 574 444 626 482
rect 574 436 583 444
rect 583 436 617 444
rect 617 436 626 444
rect 574 410 583 424
rect 583 410 617 424
rect 617 410 626 424
rect 574 372 626 410
rect 574 338 583 360
rect 583 338 617 360
rect 617 338 626 360
rect 574 308 626 338
rect 574 266 583 296
rect 583 266 617 296
rect 617 266 626 296
rect 574 244 626 266
rect 574 228 626 232
rect 574 194 583 228
rect 583 194 617 228
rect 617 194 626 228
rect 574 180 626 194
rect 574 156 626 168
rect 574 122 583 156
rect 583 122 617 156
rect 617 122 626 156
rect 574 116 626 122
<< metal2 >>
rect 10 1098 766 1104
rect 10 1046 256 1098
rect 308 1046 468 1098
rect 520 1046 766 1098
rect 10 1034 766 1046
rect 10 982 256 1034
rect 308 982 468 1034
rect 520 982 766 1034
rect 10 970 766 982
rect 10 918 256 970
rect 308 918 468 970
rect 520 918 766 970
rect 10 906 766 918
rect 10 854 256 906
rect 308 854 468 906
rect 520 854 766 906
rect 10 842 766 854
rect 10 790 256 842
rect 308 790 468 842
rect 520 790 766 842
rect 10 778 766 790
rect 10 726 256 778
rect 308 726 468 778
rect 520 726 766 778
rect 10 714 766 726
rect 10 662 256 714
rect 308 662 468 714
rect 520 662 766 714
rect 10 632 766 662
rect 10 552 766 582
rect 10 500 150 552
rect 202 500 362 552
rect 414 500 574 552
rect 626 500 766 552
rect 10 488 766 500
rect 10 436 150 488
rect 202 436 362 488
rect 414 436 574 488
rect 626 436 766 488
rect 10 424 766 436
rect 10 372 150 424
rect 202 372 362 424
rect 414 372 574 424
rect 626 372 766 424
rect 10 360 766 372
rect 10 308 150 360
rect 202 308 362 360
rect 414 308 574 360
rect 626 308 766 360
rect 10 296 766 308
rect 10 244 150 296
rect 202 244 362 296
rect 414 244 574 296
rect 626 244 766 296
rect 10 232 766 244
rect 10 180 150 232
rect 202 180 362 232
rect 414 180 574 232
rect 626 180 766 232
rect 10 168 766 180
rect 10 116 150 168
rect 202 116 362 168
rect 414 116 574 168
rect 626 116 766 168
rect 10 110 766 116
<< labels >>
flabel comment s 176 607 176 607 0 FreeSans 300 0 0 0 S
flabel comment s 176 607 176 607 0 FreeSans 300 0 0 0 S
flabel comment s 282 607 282 607 0 FreeSans 300 0 0 0 S
flabel comment s 282 607 282 607 0 FreeSans 300 0 0 0 D
flabel comment s 388 607 388 607 0 FreeSans 300 0 0 0 S
flabel comment s 388 607 388 607 0 FreeSans 300 0 0 0 S
flabel comment s 494 607 494 607 0 FreeSans 300 0 0 0 S
flabel comment s 494 607 494 607 0 FreeSans 300 0 0 0 D
flabel comment s 600 607 600 607 0 FreeSans 300 0 0 0 S
flabel metal1 s 696 603 730 614 0 FreeSans 100 0 0 0 BULK
port 2 nsew
flabel metal1 s 45 605 79 616 0 FreeSans 100 0 0 0 BULK
port 2 nsew
flabel metal1 s 368 1169 426 1194 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal1 s 349 21 407 46 0 FreeSans 100 0 0 0 GATE
port 3 nsew
flabel metal2 s 58 863 73 929 0 FreeSans 100 0 0 0 DRAIN
port 4 nsew
flabel metal2 s 51 339 65 402 0 FreeSans 100 0 0 0 SOURCE
port 5 nsew
<< properties >>
string GDS_END 9508236
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9485950
<< end >>
