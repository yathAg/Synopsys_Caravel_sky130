magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< locali >>
rect 22 992 88 1119
rect 168 1108 170 1142
rect 204 1108 266 1142
rect 300 1108 362 1142
rect 396 1108 458 1142
rect 492 1108 554 1142
rect 588 1108 650 1142
rect 684 1108 710 1142
rect 22 958 38 992
rect 72 958 88 992
rect 22 920 88 958
rect 22 886 38 920
rect 72 886 88 920
rect 22 848 88 886
rect 22 814 38 848
rect 72 814 88 848
rect 22 776 88 814
rect 22 742 38 776
rect 72 742 88 776
rect 22 704 88 742
rect 22 670 38 704
rect 72 670 88 704
rect 22 632 88 670
rect 22 598 38 632
rect 72 598 88 632
rect 22 560 88 598
rect 22 526 38 560
rect 72 526 88 560
rect 22 399 88 526
rect 792 992 858 1119
rect 792 958 808 992
rect 842 958 858 992
rect 792 920 858 958
rect 792 886 808 920
rect 842 886 858 920
rect 792 848 858 886
rect 792 814 808 848
rect 842 814 858 848
rect 792 776 858 814
rect 792 742 808 776
rect 842 742 858 776
rect 792 704 858 742
rect 792 670 808 704
rect 842 670 858 704
rect 792 632 858 670
rect 792 598 808 632
rect 842 598 858 632
rect 792 560 858 598
rect 792 526 808 560
rect 842 526 858 560
rect 168 376 170 410
rect 204 376 266 410
rect 300 376 362 410
rect 396 376 458 410
rect 492 376 554 410
rect 588 376 650 410
rect 684 376 710 410
rect 792 399 858 526
<< viali >>
rect 170 1108 204 1142
rect 266 1108 300 1142
rect 362 1108 396 1142
rect 458 1108 492 1142
rect 554 1108 588 1142
rect 650 1108 684 1142
rect 38 958 72 992
rect 38 886 72 920
rect 38 814 72 848
rect 38 742 72 776
rect 38 670 72 704
rect 38 598 72 632
rect 38 526 72 560
rect 808 958 842 992
rect 808 886 842 920
rect 808 814 842 848
rect 808 742 842 776
rect 808 670 842 704
rect 808 598 842 632
rect 808 526 842 560
rect 170 376 204 410
rect 266 376 300 410
rect 362 376 396 410
rect 458 376 492 410
rect 554 376 588 410
rect 650 376 684 410
<< obsli1 >>
rect 138 454 183 1064
rect 233 454 339 1064
rect 387 454 493 1064
rect 541 454 647 1064
rect 697 454 742 1064
<< metal1 >>
rect 164 1142 690 1154
rect 164 1108 170 1142
rect 204 1108 266 1142
rect 300 1108 362 1142
rect 396 1108 458 1142
rect 492 1108 554 1142
rect 588 1108 650 1142
rect 684 1108 690 1142
rect 164 1096 690 1108
rect 26 992 84 998
rect 26 958 38 992
rect 72 958 84 992
rect 26 920 84 958
rect 26 886 38 920
rect 72 886 84 920
rect 26 848 84 886
rect 26 814 38 848
rect 72 814 84 848
rect 26 776 84 814
rect 26 742 38 776
rect 72 742 84 776
rect 26 704 84 742
rect 26 670 38 704
rect 72 670 84 704
rect 26 632 84 670
rect 26 598 38 632
rect 72 598 84 632
rect 26 560 84 598
rect 26 526 38 560
rect 72 526 84 560
rect 26 520 84 526
rect 796 992 854 998
rect 796 958 808 992
rect 842 958 854 992
rect 796 920 854 958
rect 796 886 808 920
rect 842 886 854 920
rect 796 848 854 886
rect 796 814 808 848
rect 842 814 854 848
rect 796 776 854 814
rect 796 742 808 776
rect 842 742 854 776
rect 796 704 854 742
rect 796 670 808 704
rect 842 670 854 704
rect 796 632 854 670
rect 796 598 808 632
rect 842 598 854 632
rect 796 560 854 598
rect 796 526 808 560
rect 842 526 854 560
rect 796 520 854 526
rect 164 410 690 422
rect 164 376 170 410
rect 204 376 266 410
rect 300 376 362 410
rect 396 376 458 410
rect 492 376 554 410
rect 588 376 650 410
rect 684 376 690 410
rect 164 364 690 376
<< obsm1 >>
rect 138 722 194 1060
rect 130 466 194 722
rect 138 458 194 466
rect 223 458 349 1060
rect 377 458 503 1060
rect 531 458 657 1060
rect 686 722 742 1060
rect 686 466 750 722
rect 686 458 742 466
<< metal2 >>
rect 0 796 880 1052
rect 0 466 880 722
<< labels >>
rlabel viali s 808 958 842 992 6 BULK
port 4 nsew
rlabel viali s 808 886 842 920 6 BULK
port 4 nsew
rlabel viali s 808 814 842 848 6 BULK
port 4 nsew
rlabel viali s 808 742 842 776 6 BULK
port 4 nsew
rlabel viali s 808 670 842 704 6 BULK
port 4 nsew
rlabel viali s 808 598 842 632 6 BULK
port 4 nsew
rlabel viali s 808 526 842 560 6 BULK
port 4 nsew
rlabel viali s 38 958 72 992 6 BULK
port 4 nsew
rlabel viali s 38 886 72 920 6 BULK
port 4 nsew
rlabel viali s 38 814 72 848 6 BULK
port 4 nsew
rlabel viali s 38 742 72 776 6 BULK
port 4 nsew
rlabel viali s 38 670 72 704 6 BULK
port 4 nsew
rlabel viali s 38 598 72 632 6 BULK
port 4 nsew
rlabel viali s 38 526 72 560 6 BULK
port 4 nsew
rlabel locali s 792 399 858 1119 6 BULK
port 4 nsew
rlabel locali s 22 399 88 1119 6 BULK
port 4 nsew
rlabel metal1 s 796 520 854 998 6 BULK
port 4 nsew
rlabel metal1 s 26 520 84 998 6 BULK
port 4 nsew
rlabel metal2 s 0 796 880 1052 6 DRAIN
port 1 nsew
rlabel viali s 650 1108 684 1142 6 GATE
port 2 nsew
rlabel viali s 650 376 684 410 6 GATE
port 2 nsew
rlabel viali s 554 1108 588 1142 6 GATE
port 2 nsew
rlabel viali s 554 376 588 410 6 GATE
port 2 nsew
rlabel viali s 458 1108 492 1142 6 GATE
port 2 nsew
rlabel viali s 458 376 492 410 6 GATE
port 2 nsew
rlabel viali s 362 1108 396 1142 6 GATE
port 2 nsew
rlabel viali s 362 376 396 410 6 GATE
port 2 nsew
rlabel viali s 266 1108 300 1142 6 GATE
port 2 nsew
rlabel viali s 266 376 300 410 6 GATE
port 2 nsew
rlabel viali s 170 1108 204 1142 6 GATE
port 2 nsew
rlabel viali s 170 376 204 410 6 GATE
port 2 nsew
rlabel locali s 168 1108 710 1142 6 GATE
port 2 nsew
rlabel locali s 168 376 710 410 6 GATE
port 2 nsew
rlabel metal1 s 164 1096 690 1154 6 GATE
port 2 nsew
rlabel metal1 s 164 364 690 422 6 GATE
port 2 nsew
rlabel metal2 s 0 466 880 722 6 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX -10 0 890 1518
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10044728
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10023934
<< end >>
