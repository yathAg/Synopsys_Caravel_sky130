magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< pwell >>
rect 15 163 2283 1633
<< mvnmos >>
rect 241 189 341 1607
rect 397 189 497 1607
rect 553 189 653 1607
rect 709 189 809 1607
rect 865 189 965 1607
rect 1021 189 1121 1607
rect 1177 189 1277 1607
rect 1333 189 1433 1607
rect 1489 189 1589 1607
rect 1645 189 1745 1607
rect 1801 189 1901 1607
rect 1957 189 2057 1607
<< mvndiff >>
rect 181 1595 241 1607
rect 181 1561 196 1595
rect 230 1561 241 1595
rect 181 1527 241 1561
rect 181 1493 196 1527
rect 230 1493 241 1527
rect 181 1459 241 1493
rect 181 1425 196 1459
rect 230 1425 241 1459
rect 181 1391 241 1425
rect 181 1357 196 1391
rect 230 1357 241 1391
rect 181 1323 241 1357
rect 181 1289 196 1323
rect 230 1289 241 1323
rect 181 1255 241 1289
rect 181 1221 196 1255
rect 230 1221 241 1255
rect 181 1187 241 1221
rect 181 1153 196 1187
rect 230 1153 241 1187
rect 181 1119 241 1153
rect 181 1085 196 1119
rect 230 1085 241 1119
rect 181 1051 241 1085
rect 181 1017 196 1051
rect 230 1017 241 1051
rect 181 983 241 1017
rect 181 949 196 983
rect 230 949 241 983
rect 181 915 241 949
rect 181 881 196 915
rect 230 881 241 915
rect 181 847 241 881
rect 181 813 196 847
rect 230 813 241 847
rect 181 779 241 813
rect 181 745 196 779
rect 230 745 241 779
rect 181 711 241 745
rect 181 677 196 711
rect 230 677 241 711
rect 181 643 241 677
rect 181 609 196 643
rect 230 609 241 643
rect 181 575 241 609
rect 181 541 196 575
rect 230 541 241 575
rect 181 507 241 541
rect 181 473 196 507
rect 230 473 241 507
rect 181 439 241 473
rect 181 405 196 439
rect 230 405 241 439
rect 181 371 241 405
rect 181 337 196 371
rect 230 337 241 371
rect 181 303 241 337
rect 181 269 196 303
rect 230 269 241 303
rect 181 235 241 269
rect 181 201 196 235
rect 230 201 241 235
rect 181 189 241 201
rect 341 1595 397 1607
rect 341 1561 352 1595
rect 386 1561 397 1595
rect 341 1527 397 1561
rect 341 1493 352 1527
rect 386 1493 397 1527
rect 341 1459 397 1493
rect 341 1425 352 1459
rect 386 1425 397 1459
rect 341 1391 397 1425
rect 341 1357 352 1391
rect 386 1357 397 1391
rect 341 1323 397 1357
rect 341 1289 352 1323
rect 386 1289 397 1323
rect 341 1255 397 1289
rect 341 1221 352 1255
rect 386 1221 397 1255
rect 341 1187 397 1221
rect 341 1153 352 1187
rect 386 1153 397 1187
rect 341 1119 397 1153
rect 341 1085 352 1119
rect 386 1085 397 1119
rect 341 1051 397 1085
rect 341 1017 352 1051
rect 386 1017 397 1051
rect 341 983 397 1017
rect 341 949 352 983
rect 386 949 397 983
rect 341 915 397 949
rect 341 881 352 915
rect 386 881 397 915
rect 341 847 397 881
rect 341 813 352 847
rect 386 813 397 847
rect 341 779 397 813
rect 341 745 352 779
rect 386 745 397 779
rect 341 711 397 745
rect 341 677 352 711
rect 386 677 397 711
rect 341 643 397 677
rect 341 609 352 643
rect 386 609 397 643
rect 341 575 397 609
rect 341 541 352 575
rect 386 541 397 575
rect 341 507 397 541
rect 341 473 352 507
rect 386 473 397 507
rect 341 439 397 473
rect 341 405 352 439
rect 386 405 397 439
rect 341 371 397 405
rect 341 337 352 371
rect 386 337 397 371
rect 341 303 397 337
rect 341 269 352 303
rect 386 269 397 303
rect 341 235 397 269
rect 341 201 352 235
rect 386 201 397 235
rect 341 189 397 201
rect 497 1595 553 1607
rect 497 1561 508 1595
rect 542 1561 553 1595
rect 497 1527 553 1561
rect 497 1493 508 1527
rect 542 1493 553 1527
rect 497 1459 553 1493
rect 497 1425 508 1459
rect 542 1425 553 1459
rect 497 1391 553 1425
rect 497 1357 508 1391
rect 542 1357 553 1391
rect 497 1323 553 1357
rect 497 1289 508 1323
rect 542 1289 553 1323
rect 497 1255 553 1289
rect 497 1221 508 1255
rect 542 1221 553 1255
rect 497 1187 553 1221
rect 497 1153 508 1187
rect 542 1153 553 1187
rect 497 1119 553 1153
rect 497 1085 508 1119
rect 542 1085 553 1119
rect 497 1051 553 1085
rect 497 1017 508 1051
rect 542 1017 553 1051
rect 497 983 553 1017
rect 497 949 508 983
rect 542 949 553 983
rect 497 915 553 949
rect 497 881 508 915
rect 542 881 553 915
rect 497 847 553 881
rect 497 813 508 847
rect 542 813 553 847
rect 497 779 553 813
rect 497 745 508 779
rect 542 745 553 779
rect 497 711 553 745
rect 497 677 508 711
rect 542 677 553 711
rect 497 643 553 677
rect 497 609 508 643
rect 542 609 553 643
rect 497 575 553 609
rect 497 541 508 575
rect 542 541 553 575
rect 497 507 553 541
rect 497 473 508 507
rect 542 473 553 507
rect 497 439 553 473
rect 497 405 508 439
rect 542 405 553 439
rect 497 371 553 405
rect 497 337 508 371
rect 542 337 553 371
rect 497 303 553 337
rect 497 269 508 303
rect 542 269 553 303
rect 497 235 553 269
rect 497 201 508 235
rect 542 201 553 235
rect 497 189 553 201
rect 653 1595 709 1607
rect 653 1561 664 1595
rect 698 1561 709 1595
rect 653 1527 709 1561
rect 653 1493 664 1527
rect 698 1493 709 1527
rect 653 1459 709 1493
rect 653 1425 664 1459
rect 698 1425 709 1459
rect 653 1391 709 1425
rect 653 1357 664 1391
rect 698 1357 709 1391
rect 653 1323 709 1357
rect 653 1289 664 1323
rect 698 1289 709 1323
rect 653 1255 709 1289
rect 653 1221 664 1255
rect 698 1221 709 1255
rect 653 1187 709 1221
rect 653 1153 664 1187
rect 698 1153 709 1187
rect 653 1119 709 1153
rect 653 1085 664 1119
rect 698 1085 709 1119
rect 653 1051 709 1085
rect 653 1017 664 1051
rect 698 1017 709 1051
rect 653 983 709 1017
rect 653 949 664 983
rect 698 949 709 983
rect 653 915 709 949
rect 653 881 664 915
rect 698 881 709 915
rect 653 847 709 881
rect 653 813 664 847
rect 698 813 709 847
rect 653 779 709 813
rect 653 745 664 779
rect 698 745 709 779
rect 653 711 709 745
rect 653 677 664 711
rect 698 677 709 711
rect 653 643 709 677
rect 653 609 664 643
rect 698 609 709 643
rect 653 575 709 609
rect 653 541 664 575
rect 698 541 709 575
rect 653 507 709 541
rect 653 473 664 507
rect 698 473 709 507
rect 653 439 709 473
rect 653 405 664 439
rect 698 405 709 439
rect 653 371 709 405
rect 653 337 664 371
rect 698 337 709 371
rect 653 303 709 337
rect 653 269 664 303
rect 698 269 709 303
rect 653 235 709 269
rect 653 201 664 235
rect 698 201 709 235
rect 653 189 709 201
rect 809 1595 865 1607
rect 809 1561 820 1595
rect 854 1561 865 1595
rect 809 1527 865 1561
rect 809 1493 820 1527
rect 854 1493 865 1527
rect 809 1459 865 1493
rect 809 1425 820 1459
rect 854 1425 865 1459
rect 809 1391 865 1425
rect 809 1357 820 1391
rect 854 1357 865 1391
rect 809 1323 865 1357
rect 809 1289 820 1323
rect 854 1289 865 1323
rect 809 1255 865 1289
rect 809 1221 820 1255
rect 854 1221 865 1255
rect 809 1187 865 1221
rect 809 1153 820 1187
rect 854 1153 865 1187
rect 809 1119 865 1153
rect 809 1085 820 1119
rect 854 1085 865 1119
rect 809 1051 865 1085
rect 809 1017 820 1051
rect 854 1017 865 1051
rect 809 983 865 1017
rect 809 949 820 983
rect 854 949 865 983
rect 809 915 865 949
rect 809 881 820 915
rect 854 881 865 915
rect 809 847 865 881
rect 809 813 820 847
rect 854 813 865 847
rect 809 779 865 813
rect 809 745 820 779
rect 854 745 865 779
rect 809 711 865 745
rect 809 677 820 711
rect 854 677 865 711
rect 809 643 865 677
rect 809 609 820 643
rect 854 609 865 643
rect 809 575 865 609
rect 809 541 820 575
rect 854 541 865 575
rect 809 507 865 541
rect 809 473 820 507
rect 854 473 865 507
rect 809 439 865 473
rect 809 405 820 439
rect 854 405 865 439
rect 809 371 865 405
rect 809 337 820 371
rect 854 337 865 371
rect 809 303 865 337
rect 809 269 820 303
rect 854 269 865 303
rect 809 235 865 269
rect 809 201 820 235
rect 854 201 865 235
rect 809 189 865 201
rect 965 1595 1021 1607
rect 965 1561 976 1595
rect 1010 1561 1021 1595
rect 965 1527 1021 1561
rect 965 1493 976 1527
rect 1010 1493 1021 1527
rect 965 1459 1021 1493
rect 965 1425 976 1459
rect 1010 1425 1021 1459
rect 965 1391 1021 1425
rect 965 1357 976 1391
rect 1010 1357 1021 1391
rect 965 1323 1021 1357
rect 965 1289 976 1323
rect 1010 1289 1021 1323
rect 965 1255 1021 1289
rect 965 1221 976 1255
rect 1010 1221 1021 1255
rect 965 1187 1021 1221
rect 965 1153 976 1187
rect 1010 1153 1021 1187
rect 965 1119 1021 1153
rect 965 1085 976 1119
rect 1010 1085 1021 1119
rect 965 1051 1021 1085
rect 965 1017 976 1051
rect 1010 1017 1021 1051
rect 965 983 1021 1017
rect 965 949 976 983
rect 1010 949 1021 983
rect 965 915 1021 949
rect 965 881 976 915
rect 1010 881 1021 915
rect 965 847 1021 881
rect 965 813 976 847
rect 1010 813 1021 847
rect 965 779 1021 813
rect 965 745 976 779
rect 1010 745 1021 779
rect 965 711 1021 745
rect 965 677 976 711
rect 1010 677 1021 711
rect 965 643 1021 677
rect 965 609 976 643
rect 1010 609 1021 643
rect 965 575 1021 609
rect 965 541 976 575
rect 1010 541 1021 575
rect 965 507 1021 541
rect 965 473 976 507
rect 1010 473 1021 507
rect 965 439 1021 473
rect 965 405 976 439
rect 1010 405 1021 439
rect 965 371 1021 405
rect 965 337 976 371
rect 1010 337 1021 371
rect 965 303 1021 337
rect 965 269 976 303
rect 1010 269 1021 303
rect 965 235 1021 269
rect 965 201 976 235
rect 1010 201 1021 235
rect 965 189 1021 201
rect 1121 1595 1177 1607
rect 1121 1561 1132 1595
rect 1166 1561 1177 1595
rect 1121 1527 1177 1561
rect 1121 1493 1132 1527
rect 1166 1493 1177 1527
rect 1121 1459 1177 1493
rect 1121 1425 1132 1459
rect 1166 1425 1177 1459
rect 1121 1391 1177 1425
rect 1121 1357 1132 1391
rect 1166 1357 1177 1391
rect 1121 1323 1177 1357
rect 1121 1289 1132 1323
rect 1166 1289 1177 1323
rect 1121 1255 1177 1289
rect 1121 1221 1132 1255
rect 1166 1221 1177 1255
rect 1121 1187 1177 1221
rect 1121 1153 1132 1187
rect 1166 1153 1177 1187
rect 1121 1119 1177 1153
rect 1121 1085 1132 1119
rect 1166 1085 1177 1119
rect 1121 1051 1177 1085
rect 1121 1017 1132 1051
rect 1166 1017 1177 1051
rect 1121 983 1177 1017
rect 1121 949 1132 983
rect 1166 949 1177 983
rect 1121 915 1177 949
rect 1121 881 1132 915
rect 1166 881 1177 915
rect 1121 847 1177 881
rect 1121 813 1132 847
rect 1166 813 1177 847
rect 1121 779 1177 813
rect 1121 745 1132 779
rect 1166 745 1177 779
rect 1121 711 1177 745
rect 1121 677 1132 711
rect 1166 677 1177 711
rect 1121 643 1177 677
rect 1121 609 1132 643
rect 1166 609 1177 643
rect 1121 575 1177 609
rect 1121 541 1132 575
rect 1166 541 1177 575
rect 1121 507 1177 541
rect 1121 473 1132 507
rect 1166 473 1177 507
rect 1121 439 1177 473
rect 1121 405 1132 439
rect 1166 405 1177 439
rect 1121 371 1177 405
rect 1121 337 1132 371
rect 1166 337 1177 371
rect 1121 303 1177 337
rect 1121 269 1132 303
rect 1166 269 1177 303
rect 1121 235 1177 269
rect 1121 201 1132 235
rect 1166 201 1177 235
rect 1121 189 1177 201
rect 1277 1595 1333 1607
rect 1277 1561 1288 1595
rect 1322 1561 1333 1595
rect 1277 1527 1333 1561
rect 1277 1493 1288 1527
rect 1322 1493 1333 1527
rect 1277 1459 1333 1493
rect 1277 1425 1288 1459
rect 1322 1425 1333 1459
rect 1277 1391 1333 1425
rect 1277 1357 1288 1391
rect 1322 1357 1333 1391
rect 1277 1323 1333 1357
rect 1277 1289 1288 1323
rect 1322 1289 1333 1323
rect 1277 1255 1333 1289
rect 1277 1221 1288 1255
rect 1322 1221 1333 1255
rect 1277 1187 1333 1221
rect 1277 1153 1288 1187
rect 1322 1153 1333 1187
rect 1277 1119 1333 1153
rect 1277 1085 1288 1119
rect 1322 1085 1333 1119
rect 1277 1051 1333 1085
rect 1277 1017 1288 1051
rect 1322 1017 1333 1051
rect 1277 983 1333 1017
rect 1277 949 1288 983
rect 1322 949 1333 983
rect 1277 915 1333 949
rect 1277 881 1288 915
rect 1322 881 1333 915
rect 1277 847 1333 881
rect 1277 813 1288 847
rect 1322 813 1333 847
rect 1277 779 1333 813
rect 1277 745 1288 779
rect 1322 745 1333 779
rect 1277 711 1333 745
rect 1277 677 1288 711
rect 1322 677 1333 711
rect 1277 643 1333 677
rect 1277 609 1288 643
rect 1322 609 1333 643
rect 1277 575 1333 609
rect 1277 541 1288 575
rect 1322 541 1333 575
rect 1277 507 1333 541
rect 1277 473 1288 507
rect 1322 473 1333 507
rect 1277 439 1333 473
rect 1277 405 1288 439
rect 1322 405 1333 439
rect 1277 371 1333 405
rect 1277 337 1288 371
rect 1322 337 1333 371
rect 1277 303 1333 337
rect 1277 269 1288 303
rect 1322 269 1333 303
rect 1277 235 1333 269
rect 1277 201 1288 235
rect 1322 201 1333 235
rect 1277 189 1333 201
rect 1433 1595 1489 1607
rect 1433 1561 1444 1595
rect 1478 1561 1489 1595
rect 1433 1527 1489 1561
rect 1433 1493 1444 1527
rect 1478 1493 1489 1527
rect 1433 1459 1489 1493
rect 1433 1425 1444 1459
rect 1478 1425 1489 1459
rect 1433 1391 1489 1425
rect 1433 1357 1444 1391
rect 1478 1357 1489 1391
rect 1433 1323 1489 1357
rect 1433 1289 1444 1323
rect 1478 1289 1489 1323
rect 1433 1255 1489 1289
rect 1433 1221 1444 1255
rect 1478 1221 1489 1255
rect 1433 1187 1489 1221
rect 1433 1153 1444 1187
rect 1478 1153 1489 1187
rect 1433 1119 1489 1153
rect 1433 1085 1444 1119
rect 1478 1085 1489 1119
rect 1433 1051 1489 1085
rect 1433 1017 1444 1051
rect 1478 1017 1489 1051
rect 1433 983 1489 1017
rect 1433 949 1444 983
rect 1478 949 1489 983
rect 1433 915 1489 949
rect 1433 881 1444 915
rect 1478 881 1489 915
rect 1433 847 1489 881
rect 1433 813 1444 847
rect 1478 813 1489 847
rect 1433 779 1489 813
rect 1433 745 1444 779
rect 1478 745 1489 779
rect 1433 711 1489 745
rect 1433 677 1444 711
rect 1478 677 1489 711
rect 1433 643 1489 677
rect 1433 609 1444 643
rect 1478 609 1489 643
rect 1433 575 1489 609
rect 1433 541 1444 575
rect 1478 541 1489 575
rect 1433 507 1489 541
rect 1433 473 1444 507
rect 1478 473 1489 507
rect 1433 439 1489 473
rect 1433 405 1444 439
rect 1478 405 1489 439
rect 1433 371 1489 405
rect 1433 337 1444 371
rect 1478 337 1489 371
rect 1433 303 1489 337
rect 1433 269 1444 303
rect 1478 269 1489 303
rect 1433 235 1489 269
rect 1433 201 1444 235
rect 1478 201 1489 235
rect 1433 189 1489 201
rect 1589 1595 1645 1607
rect 1589 1561 1600 1595
rect 1634 1561 1645 1595
rect 1589 1527 1645 1561
rect 1589 1493 1600 1527
rect 1634 1493 1645 1527
rect 1589 1459 1645 1493
rect 1589 1425 1600 1459
rect 1634 1425 1645 1459
rect 1589 1391 1645 1425
rect 1589 1357 1600 1391
rect 1634 1357 1645 1391
rect 1589 1323 1645 1357
rect 1589 1289 1600 1323
rect 1634 1289 1645 1323
rect 1589 1255 1645 1289
rect 1589 1221 1600 1255
rect 1634 1221 1645 1255
rect 1589 1187 1645 1221
rect 1589 1153 1600 1187
rect 1634 1153 1645 1187
rect 1589 1119 1645 1153
rect 1589 1085 1600 1119
rect 1634 1085 1645 1119
rect 1589 1051 1645 1085
rect 1589 1017 1600 1051
rect 1634 1017 1645 1051
rect 1589 983 1645 1017
rect 1589 949 1600 983
rect 1634 949 1645 983
rect 1589 915 1645 949
rect 1589 881 1600 915
rect 1634 881 1645 915
rect 1589 847 1645 881
rect 1589 813 1600 847
rect 1634 813 1645 847
rect 1589 779 1645 813
rect 1589 745 1600 779
rect 1634 745 1645 779
rect 1589 711 1645 745
rect 1589 677 1600 711
rect 1634 677 1645 711
rect 1589 643 1645 677
rect 1589 609 1600 643
rect 1634 609 1645 643
rect 1589 575 1645 609
rect 1589 541 1600 575
rect 1634 541 1645 575
rect 1589 507 1645 541
rect 1589 473 1600 507
rect 1634 473 1645 507
rect 1589 439 1645 473
rect 1589 405 1600 439
rect 1634 405 1645 439
rect 1589 371 1645 405
rect 1589 337 1600 371
rect 1634 337 1645 371
rect 1589 303 1645 337
rect 1589 269 1600 303
rect 1634 269 1645 303
rect 1589 235 1645 269
rect 1589 201 1600 235
rect 1634 201 1645 235
rect 1589 189 1645 201
rect 1745 1595 1801 1607
rect 1745 1561 1756 1595
rect 1790 1561 1801 1595
rect 1745 1527 1801 1561
rect 1745 1493 1756 1527
rect 1790 1493 1801 1527
rect 1745 1459 1801 1493
rect 1745 1425 1756 1459
rect 1790 1425 1801 1459
rect 1745 1391 1801 1425
rect 1745 1357 1756 1391
rect 1790 1357 1801 1391
rect 1745 1323 1801 1357
rect 1745 1289 1756 1323
rect 1790 1289 1801 1323
rect 1745 1255 1801 1289
rect 1745 1221 1756 1255
rect 1790 1221 1801 1255
rect 1745 1187 1801 1221
rect 1745 1153 1756 1187
rect 1790 1153 1801 1187
rect 1745 1119 1801 1153
rect 1745 1085 1756 1119
rect 1790 1085 1801 1119
rect 1745 1051 1801 1085
rect 1745 1017 1756 1051
rect 1790 1017 1801 1051
rect 1745 983 1801 1017
rect 1745 949 1756 983
rect 1790 949 1801 983
rect 1745 915 1801 949
rect 1745 881 1756 915
rect 1790 881 1801 915
rect 1745 847 1801 881
rect 1745 813 1756 847
rect 1790 813 1801 847
rect 1745 779 1801 813
rect 1745 745 1756 779
rect 1790 745 1801 779
rect 1745 711 1801 745
rect 1745 677 1756 711
rect 1790 677 1801 711
rect 1745 643 1801 677
rect 1745 609 1756 643
rect 1790 609 1801 643
rect 1745 575 1801 609
rect 1745 541 1756 575
rect 1790 541 1801 575
rect 1745 507 1801 541
rect 1745 473 1756 507
rect 1790 473 1801 507
rect 1745 439 1801 473
rect 1745 405 1756 439
rect 1790 405 1801 439
rect 1745 371 1801 405
rect 1745 337 1756 371
rect 1790 337 1801 371
rect 1745 303 1801 337
rect 1745 269 1756 303
rect 1790 269 1801 303
rect 1745 235 1801 269
rect 1745 201 1756 235
rect 1790 201 1801 235
rect 1745 189 1801 201
rect 1901 1595 1957 1607
rect 1901 1561 1912 1595
rect 1946 1561 1957 1595
rect 1901 1527 1957 1561
rect 1901 1493 1912 1527
rect 1946 1493 1957 1527
rect 1901 1459 1957 1493
rect 1901 1425 1912 1459
rect 1946 1425 1957 1459
rect 1901 1391 1957 1425
rect 1901 1357 1912 1391
rect 1946 1357 1957 1391
rect 1901 1323 1957 1357
rect 1901 1289 1912 1323
rect 1946 1289 1957 1323
rect 1901 1255 1957 1289
rect 1901 1221 1912 1255
rect 1946 1221 1957 1255
rect 1901 1187 1957 1221
rect 1901 1153 1912 1187
rect 1946 1153 1957 1187
rect 1901 1119 1957 1153
rect 1901 1085 1912 1119
rect 1946 1085 1957 1119
rect 1901 1051 1957 1085
rect 1901 1017 1912 1051
rect 1946 1017 1957 1051
rect 1901 983 1957 1017
rect 1901 949 1912 983
rect 1946 949 1957 983
rect 1901 915 1957 949
rect 1901 881 1912 915
rect 1946 881 1957 915
rect 1901 847 1957 881
rect 1901 813 1912 847
rect 1946 813 1957 847
rect 1901 779 1957 813
rect 1901 745 1912 779
rect 1946 745 1957 779
rect 1901 711 1957 745
rect 1901 677 1912 711
rect 1946 677 1957 711
rect 1901 643 1957 677
rect 1901 609 1912 643
rect 1946 609 1957 643
rect 1901 575 1957 609
rect 1901 541 1912 575
rect 1946 541 1957 575
rect 1901 507 1957 541
rect 1901 473 1912 507
rect 1946 473 1957 507
rect 1901 439 1957 473
rect 1901 405 1912 439
rect 1946 405 1957 439
rect 1901 371 1957 405
rect 1901 337 1912 371
rect 1946 337 1957 371
rect 1901 303 1957 337
rect 1901 269 1912 303
rect 1946 269 1957 303
rect 1901 235 1957 269
rect 1901 201 1912 235
rect 1946 201 1957 235
rect 1901 189 1957 201
rect 2057 1595 2117 1607
rect 2057 1561 2068 1595
rect 2102 1561 2117 1595
rect 2057 1527 2117 1561
rect 2057 1493 2068 1527
rect 2102 1493 2117 1527
rect 2057 1459 2117 1493
rect 2057 1425 2068 1459
rect 2102 1425 2117 1459
rect 2057 1391 2117 1425
rect 2057 1357 2068 1391
rect 2102 1357 2117 1391
rect 2057 1323 2117 1357
rect 2057 1289 2068 1323
rect 2102 1289 2117 1323
rect 2057 1255 2117 1289
rect 2057 1221 2068 1255
rect 2102 1221 2117 1255
rect 2057 1187 2117 1221
rect 2057 1153 2068 1187
rect 2102 1153 2117 1187
rect 2057 1119 2117 1153
rect 2057 1085 2068 1119
rect 2102 1085 2117 1119
rect 2057 1051 2117 1085
rect 2057 1017 2068 1051
rect 2102 1017 2117 1051
rect 2057 983 2117 1017
rect 2057 949 2068 983
rect 2102 949 2117 983
rect 2057 915 2117 949
rect 2057 881 2068 915
rect 2102 881 2117 915
rect 2057 847 2117 881
rect 2057 813 2068 847
rect 2102 813 2117 847
rect 2057 779 2117 813
rect 2057 745 2068 779
rect 2102 745 2117 779
rect 2057 711 2117 745
rect 2057 677 2068 711
rect 2102 677 2117 711
rect 2057 643 2117 677
rect 2057 609 2068 643
rect 2102 609 2117 643
rect 2057 575 2117 609
rect 2057 541 2068 575
rect 2102 541 2117 575
rect 2057 507 2117 541
rect 2057 473 2068 507
rect 2102 473 2117 507
rect 2057 439 2117 473
rect 2057 405 2068 439
rect 2102 405 2117 439
rect 2057 371 2117 405
rect 2057 337 2068 371
rect 2102 337 2117 371
rect 2057 303 2117 337
rect 2057 269 2068 303
rect 2102 269 2117 303
rect 2057 235 2117 269
rect 2057 201 2068 235
rect 2102 201 2117 235
rect 2057 189 2117 201
<< mvndiffc >>
rect 196 1561 230 1595
rect 196 1493 230 1527
rect 196 1425 230 1459
rect 196 1357 230 1391
rect 196 1289 230 1323
rect 196 1221 230 1255
rect 196 1153 230 1187
rect 196 1085 230 1119
rect 196 1017 230 1051
rect 196 949 230 983
rect 196 881 230 915
rect 196 813 230 847
rect 196 745 230 779
rect 196 677 230 711
rect 196 609 230 643
rect 196 541 230 575
rect 196 473 230 507
rect 196 405 230 439
rect 196 337 230 371
rect 196 269 230 303
rect 196 201 230 235
rect 352 1561 386 1595
rect 352 1493 386 1527
rect 352 1425 386 1459
rect 352 1357 386 1391
rect 352 1289 386 1323
rect 352 1221 386 1255
rect 352 1153 386 1187
rect 352 1085 386 1119
rect 352 1017 386 1051
rect 352 949 386 983
rect 352 881 386 915
rect 352 813 386 847
rect 352 745 386 779
rect 352 677 386 711
rect 352 609 386 643
rect 352 541 386 575
rect 352 473 386 507
rect 352 405 386 439
rect 352 337 386 371
rect 352 269 386 303
rect 352 201 386 235
rect 508 1561 542 1595
rect 508 1493 542 1527
rect 508 1425 542 1459
rect 508 1357 542 1391
rect 508 1289 542 1323
rect 508 1221 542 1255
rect 508 1153 542 1187
rect 508 1085 542 1119
rect 508 1017 542 1051
rect 508 949 542 983
rect 508 881 542 915
rect 508 813 542 847
rect 508 745 542 779
rect 508 677 542 711
rect 508 609 542 643
rect 508 541 542 575
rect 508 473 542 507
rect 508 405 542 439
rect 508 337 542 371
rect 508 269 542 303
rect 508 201 542 235
rect 664 1561 698 1595
rect 664 1493 698 1527
rect 664 1425 698 1459
rect 664 1357 698 1391
rect 664 1289 698 1323
rect 664 1221 698 1255
rect 664 1153 698 1187
rect 664 1085 698 1119
rect 664 1017 698 1051
rect 664 949 698 983
rect 664 881 698 915
rect 664 813 698 847
rect 664 745 698 779
rect 664 677 698 711
rect 664 609 698 643
rect 664 541 698 575
rect 664 473 698 507
rect 664 405 698 439
rect 664 337 698 371
rect 664 269 698 303
rect 664 201 698 235
rect 820 1561 854 1595
rect 820 1493 854 1527
rect 820 1425 854 1459
rect 820 1357 854 1391
rect 820 1289 854 1323
rect 820 1221 854 1255
rect 820 1153 854 1187
rect 820 1085 854 1119
rect 820 1017 854 1051
rect 820 949 854 983
rect 820 881 854 915
rect 820 813 854 847
rect 820 745 854 779
rect 820 677 854 711
rect 820 609 854 643
rect 820 541 854 575
rect 820 473 854 507
rect 820 405 854 439
rect 820 337 854 371
rect 820 269 854 303
rect 820 201 854 235
rect 976 1561 1010 1595
rect 976 1493 1010 1527
rect 976 1425 1010 1459
rect 976 1357 1010 1391
rect 976 1289 1010 1323
rect 976 1221 1010 1255
rect 976 1153 1010 1187
rect 976 1085 1010 1119
rect 976 1017 1010 1051
rect 976 949 1010 983
rect 976 881 1010 915
rect 976 813 1010 847
rect 976 745 1010 779
rect 976 677 1010 711
rect 976 609 1010 643
rect 976 541 1010 575
rect 976 473 1010 507
rect 976 405 1010 439
rect 976 337 1010 371
rect 976 269 1010 303
rect 976 201 1010 235
rect 1132 1561 1166 1595
rect 1132 1493 1166 1527
rect 1132 1425 1166 1459
rect 1132 1357 1166 1391
rect 1132 1289 1166 1323
rect 1132 1221 1166 1255
rect 1132 1153 1166 1187
rect 1132 1085 1166 1119
rect 1132 1017 1166 1051
rect 1132 949 1166 983
rect 1132 881 1166 915
rect 1132 813 1166 847
rect 1132 745 1166 779
rect 1132 677 1166 711
rect 1132 609 1166 643
rect 1132 541 1166 575
rect 1132 473 1166 507
rect 1132 405 1166 439
rect 1132 337 1166 371
rect 1132 269 1166 303
rect 1132 201 1166 235
rect 1288 1561 1322 1595
rect 1288 1493 1322 1527
rect 1288 1425 1322 1459
rect 1288 1357 1322 1391
rect 1288 1289 1322 1323
rect 1288 1221 1322 1255
rect 1288 1153 1322 1187
rect 1288 1085 1322 1119
rect 1288 1017 1322 1051
rect 1288 949 1322 983
rect 1288 881 1322 915
rect 1288 813 1322 847
rect 1288 745 1322 779
rect 1288 677 1322 711
rect 1288 609 1322 643
rect 1288 541 1322 575
rect 1288 473 1322 507
rect 1288 405 1322 439
rect 1288 337 1322 371
rect 1288 269 1322 303
rect 1288 201 1322 235
rect 1444 1561 1478 1595
rect 1444 1493 1478 1527
rect 1444 1425 1478 1459
rect 1444 1357 1478 1391
rect 1444 1289 1478 1323
rect 1444 1221 1478 1255
rect 1444 1153 1478 1187
rect 1444 1085 1478 1119
rect 1444 1017 1478 1051
rect 1444 949 1478 983
rect 1444 881 1478 915
rect 1444 813 1478 847
rect 1444 745 1478 779
rect 1444 677 1478 711
rect 1444 609 1478 643
rect 1444 541 1478 575
rect 1444 473 1478 507
rect 1444 405 1478 439
rect 1444 337 1478 371
rect 1444 269 1478 303
rect 1444 201 1478 235
rect 1600 1561 1634 1595
rect 1600 1493 1634 1527
rect 1600 1425 1634 1459
rect 1600 1357 1634 1391
rect 1600 1289 1634 1323
rect 1600 1221 1634 1255
rect 1600 1153 1634 1187
rect 1600 1085 1634 1119
rect 1600 1017 1634 1051
rect 1600 949 1634 983
rect 1600 881 1634 915
rect 1600 813 1634 847
rect 1600 745 1634 779
rect 1600 677 1634 711
rect 1600 609 1634 643
rect 1600 541 1634 575
rect 1600 473 1634 507
rect 1600 405 1634 439
rect 1600 337 1634 371
rect 1600 269 1634 303
rect 1600 201 1634 235
rect 1756 1561 1790 1595
rect 1756 1493 1790 1527
rect 1756 1425 1790 1459
rect 1756 1357 1790 1391
rect 1756 1289 1790 1323
rect 1756 1221 1790 1255
rect 1756 1153 1790 1187
rect 1756 1085 1790 1119
rect 1756 1017 1790 1051
rect 1756 949 1790 983
rect 1756 881 1790 915
rect 1756 813 1790 847
rect 1756 745 1790 779
rect 1756 677 1790 711
rect 1756 609 1790 643
rect 1756 541 1790 575
rect 1756 473 1790 507
rect 1756 405 1790 439
rect 1756 337 1790 371
rect 1756 269 1790 303
rect 1756 201 1790 235
rect 1912 1561 1946 1595
rect 1912 1493 1946 1527
rect 1912 1425 1946 1459
rect 1912 1357 1946 1391
rect 1912 1289 1946 1323
rect 1912 1221 1946 1255
rect 1912 1153 1946 1187
rect 1912 1085 1946 1119
rect 1912 1017 1946 1051
rect 1912 949 1946 983
rect 1912 881 1946 915
rect 1912 813 1946 847
rect 1912 745 1946 779
rect 1912 677 1946 711
rect 1912 609 1946 643
rect 1912 541 1946 575
rect 1912 473 1946 507
rect 1912 405 1946 439
rect 1912 337 1946 371
rect 1912 269 1946 303
rect 1912 201 1946 235
rect 2068 1561 2102 1595
rect 2068 1493 2102 1527
rect 2068 1425 2102 1459
rect 2068 1357 2102 1391
rect 2068 1289 2102 1323
rect 2068 1221 2102 1255
rect 2068 1153 2102 1187
rect 2068 1085 2102 1119
rect 2068 1017 2102 1051
rect 2068 949 2102 983
rect 2068 881 2102 915
rect 2068 813 2102 847
rect 2068 745 2102 779
rect 2068 677 2102 711
rect 2068 609 2102 643
rect 2068 541 2102 575
rect 2068 473 2102 507
rect 2068 405 2102 439
rect 2068 337 2102 371
rect 2068 269 2102 303
rect 2068 201 2102 235
<< mvpsubdiff >>
rect 41 1595 181 1607
rect 41 201 60 1595
rect 162 201 181 1595
rect 41 189 181 201
rect 2117 1595 2257 1607
rect 2117 201 2136 1595
rect 2238 201 2257 1595
rect 2117 189 2257 201
<< mvpsubdiffcont >>
rect 60 201 162 1595
rect 2136 201 2238 1595
<< poly >>
rect 383 1775 1915 1796
rect 190 1683 341 1699
rect 190 1649 206 1683
rect 240 1649 341 1683
rect 383 1673 418 1775
rect 1880 1673 1915 1775
rect 383 1657 1915 1673
rect 1957 1683 2108 1699
rect 190 1633 341 1649
rect 241 1607 341 1633
rect 397 1607 497 1657
rect 553 1607 653 1657
rect 709 1607 809 1657
rect 865 1607 965 1657
rect 1021 1607 1121 1657
rect 1177 1607 1277 1657
rect 1333 1607 1433 1657
rect 1489 1607 1589 1657
rect 1645 1607 1745 1657
rect 1801 1607 1901 1657
rect 1957 1649 2058 1683
rect 2092 1649 2108 1683
rect 1957 1633 2108 1649
rect 1957 1607 2057 1633
rect 241 163 341 189
rect 190 147 341 163
rect 190 113 206 147
rect 240 113 341 147
rect 397 139 497 189
rect 553 139 653 189
rect 709 139 809 189
rect 865 139 965 189
rect 1021 139 1121 189
rect 1177 139 1277 189
rect 1333 139 1433 189
rect 1489 139 1589 189
rect 1645 139 1745 189
rect 1801 139 1901 189
rect 1957 163 2057 189
rect 1957 147 2108 163
rect 190 97 341 113
rect 383 123 1915 139
rect 383 21 418 123
rect 1880 21 1915 123
rect 1957 113 2058 147
rect 2092 113 2108 147
rect 1957 97 2108 113
rect 383 0 1915 21
<< polycont >>
rect 206 1649 240 1683
rect 418 1673 1880 1775
rect 2058 1649 2092 1683
rect 206 113 240 147
rect 418 21 1880 123
rect 2058 113 2092 147
<< locali >>
rect 385 1777 1913 1796
rect 190 1683 256 1699
rect 190 1649 206 1683
rect 240 1649 256 1683
rect 385 1671 412 1777
rect 1886 1671 1913 1777
rect 385 1659 1913 1671
rect 2042 1683 2108 1699
rect 190 1633 256 1649
rect 2042 1649 2058 1683
rect 2092 1649 2108 1683
rect 2042 1633 2108 1649
rect 190 1611 230 1633
rect 2068 1611 2108 1633
rect 41 1595 230 1611
rect 41 201 60 1595
rect 162 1561 196 1595
rect 162 1527 230 1561
rect 162 1493 196 1527
rect 162 1459 230 1493
rect 162 1425 196 1459
rect 162 1391 230 1425
rect 162 1357 196 1391
rect 162 1323 230 1357
rect 162 1289 196 1323
rect 162 1255 230 1289
rect 162 1221 196 1255
rect 162 1187 230 1221
rect 162 1153 196 1187
rect 162 1119 230 1153
rect 162 1085 196 1119
rect 162 1051 230 1085
rect 162 1017 196 1051
rect 162 983 230 1017
rect 162 949 196 983
rect 162 915 230 949
rect 162 881 196 915
rect 162 847 230 881
rect 162 813 196 847
rect 162 779 230 813
rect 162 745 196 779
rect 162 711 230 745
rect 162 677 196 711
rect 162 643 230 677
rect 162 609 196 643
rect 162 575 230 609
rect 162 541 196 575
rect 162 507 230 541
rect 162 473 196 507
rect 162 439 230 473
rect 162 405 196 439
rect 162 371 230 405
rect 162 337 196 371
rect 162 303 230 337
rect 162 269 196 303
rect 162 235 230 269
rect 162 201 196 235
rect 41 185 230 201
rect 352 1595 386 1611
rect 352 1527 386 1529
rect 352 1491 386 1493
rect 352 1419 386 1425
rect 352 1347 386 1357
rect 352 1275 386 1289
rect 352 1203 386 1221
rect 352 1131 386 1153
rect 352 1059 386 1085
rect 352 987 386 1017
rect 352 915 386 949
rect 352 847 386 881
rect 352 779 386 809
rect 352 711 386 737
rect 352 643 386 665
rect 352 575 386 593
rect 352 507 386 521
rect 352 439 386 449
rect 352 371 386 377
rect 352 303 386 305
rect 352 267 386 269
rect 352 185 386 201
rect 508 1595 542 1611
rect 508 1527 542 1529
rect 508 1491 542 1493
rect 508 1419 542 1425
rect 508 1347 542 1357
rect 508 1275 542 1289
rect 508 1203 542 1221
rect 508 1131 542 1153
rect 508 1059 542 1085
rect 508 987 542 1017
rect 508 915 542 949
rect 508 847 542 881
rect 508 779 542 809
rect 508 711 542 737
rect 508 643 542 665
rect 508 575 542 593
rect 508 507 542 521
rect 508 439 542 449
rect 508 371 542 377
rect 508 303 542 305
rect 508 267 542 269
rect 508 185 542 201
rect 664 1595 698 1611
rect 664 1527 698 1529
rect 664 1491 698 1493
rect 664 1419 698 1425
rect 664 1347 698 1357
rect 664 1275 698 1289
rect 664 1203 698 1221
rect 664 1131 698 1153
rect 664 1059 698 1085
rect 664 987 698 1017
rect 664 915 698 949
rect 664 847 698 881
rect 664 779 698 809
rect 664 711 698 737
rect 664 643 698 665
rect 664 575 698 593
rect 664 507 698 521
rect 664 439 698 449
rect 664 371 698 377
rect 664 303 698 305
rect 664 267 698 269
rect 664 185 698 201
rect 820 1595 854 1611
rect 820 1527 854 1529
rect 820 1491 854 1493
rect 820 1419 854 1425
rect 820 1347 854 1357
rect 820 1275 854 1289
rect 820 1203 854 1221
rect 820 1131 854 1153
rect 820 1059 854 1085
rect 820 987 854 1017
rect 820 915 854 949
rect 820 847 854 881
rect 820 779 854 809
rect 820 711 854 737
rect 820 643 854 665
rect 820 575 854 593
rect 820 507 854 521
rect 820 439 854 449
rect 820 371 854 377
rect 820 303 854 305
rect 820 267 854 269
rect 820 185 854 201
rect 976 1595 1010 1611
rect 976 1527 1010 1529
rect 976 1491 1010 1493
rect 976 1419 1010 1425
rect 976 1347 1010 1357
rect 976 1275 1010 1289
rect 976 1203 1010 1221
rect 976 1131 1010 1153
rect 976 1059 1010 1085
rect 976 987 1010 1017
rect 976 915 1010 949
rect 976 847 1010 881
rect 976 779 1010 809
rect 976 711 1010 737
rect 976 643 1010 665
rect 976 575 1010 593
rect 976 507 1010 521
rect 976 439 1010 449
rect 976 371 1010 377
rect 976 303 1010 305
rect 976 267 1010 269
rect 976 185 1010 201
rect 1132 1595 1166 1611
rect 1132 1527 1166 1529
rect 1132 1491 1166 1493
rect 1132 1419 1166 1425
rect 1132 1347 1166 1357
rect 1132 1275 1166 1289
rect 1132 1203 1166 1221
rect 1132 1131 1166 1153
rect 1132 1059 1166 1085
rect 1132 987 1166 1017
rect 1132 915 1166 949
rect 1132 847 1166 881
rect 1132 779 1166 809
rect 1132 711 1166 737
rect 1132 643 1166 665
rect 1132 575 1166 593
rect 1132 507 1166 521
rect 1132 439 1166 449
rect 1132 371 1166 377
rect 1132 303 1166 305
rect 1132 267 1166 269
rect 1132 185 1166 201
rect 1288 1595 1322 1611
rect 1288 1527 1322 1529
rect 1288 1491 1322 1493
rect 1288 1419 1322 1425
rect 1288 1347 1322 1357
rect 1288 1275 1322 1289
rect 1288 1203 1322 1221
rect 1288 1131 1322 1153
rect 1288 1059 1322 1085
rect 1288 987 1322 1017
rect 1288 915 1322 949
rect 1288 847 1322 881
rect 1288 779 1322 809
rect 1288 711 1322 737
rect 1288 643 1322 665
rect 1288 575 1322 593
rect 1288 507 1322 521
rect 1288 439 1322 449
rect 1288 371 1322 377
rect 1288 303 1322 305
rect 1288 267 1322 269
rect 1288 185 1322 201
rect 1444 1595 1478 1611
rect 1444 1527 1478 1529
rect 1444 1491 1478 1493
rect 1444 1419 1478 1425
rect 1444 1347 1478 1357
rect 1444 1275 1478 1289
rect 1444 1203 1478 1221
rect 1444 1131 1478 1153
rect 1444 1059 1478 1085
rect 1444 987 1478 1017
rect 1444 915 1478 949
rect 1444 847 1478 881
rect 1444 779 1478 809
rect 1444 711 1478 737
rect 1444 643 1478 665
rect 1444 575 1478 593
rect 1444 507 1478 521
rect 1444 439 1478 449
rect 1444 371 1478 377
rect 1444 303 1478 305
rect 1444 267 1478 269
rect 1444 185 1478 201
rect 1600 1595 1634 1611
rect 1600 1527 1634 1529
rect 1600 1491 1634 1493
rect 1600 1419 1634 1425
rect 1600 1347 1634 1357
rect 1600 1275 1634 1289
rect 1600 1203 1634 1221
rect 1600 1131 1634 1153
rect 1600 1059 1634 1085
rect 1600 987 1634 1017
rect 1600 915 1634 949
rect 1600 847 1634 881
rect 1600 779 1634 809
rect 1600 711 1634 737
rect 1600 643 1634 665
rect 1600 575 1634 593
rect 1600 507 1634 521
rect 1600 439 1634 449
rect 1600 371 1634 377
rect 1600 303 1634 305
rect 1600 267 1634 269
rect 1600 185 1634 201
rect 1756 1595 1790 1611
rect 1756 1527 1790 1529
rect 1756 1491 1790 1493
rect 1756 1419 1790 1425
rect 1756 1347 1790 1357
rect 1756 1275 1790 1289
rect 1756 1203 1790 1221
rect 1756 1131 1790 1153
rect 1756 1059 1790 1085
rect 1756 987 1790 1017
rect 1756 915 1790 949
rect 1756 847 1790 881
rect 1756 779 1790 809
rect 1756 711 1790 737
rect 1756 643 1790 665
rect 1756 575 1790 593
rect 1756 507 1790 521
rect 1756 439 1790 449
rect 1756 371 1790 377
rect 1756 303 1790 305
rect 1756 267 1790 269
rect 1756 185 1790 201
rect 1912 1595 1946 1611
rect 1912 1527 1946 1529
rect 1912 1491 1946 1493
rect 1912 1419 1946 1425
rect 1912 1347 1946 1357
rect 1912 1275 1946 1289
rect 1912 1203 1946 1221
rect 1912 1131 1946 1153
rect 1912 1059 1946 1085
rect 1912 987 1946 1017
rect 1912 915 1946 949
rect 1912 847 1946 881
rect 1912 779 1946 809
rect 1912 711 1946 737
rect 1912 643 1946 665
rect 1912 575 1946 593
rect 1912 507 1946 521
rect 1912 439 1946 449
rect 1912 371 1946 377
rect 1912 303 1946 305
rect 1912 267 1946 269
rect 1912 185 1946 201
rect 2068 1595 2257 1611
rect 2102 1561 2136 1595
rect 2068 1527 2136 1561
rect 2102 1493 2136 1527
rect 2068 1459 2136 1493
rect 2102 1425 2136 1459
rect 2068 1391 2136 1425
rect 2102 1357 2136 1391
rect 2068 1323 2136 1357
rect 2102 1289 2136 1323
rect 2068 1255 2136 1289
rect 2102 1221 2136 1255
rect 2068 1187 2136 1221
rect 2102 1153 2136 1187
rect 2068 1119 2136 1153
rect 2102 1085 2136 1119
rect 2068 1051 2136 1085
rect 2102 1017 2136 1051
rect 2068 983 2136 1017
rect 2102 949 2136 983
rect 2068 915 2136 949
rect 2102 881 2136 915
rect 2068 847 2136 881
rect 2102 813 2136 847
rect 2068 779 2136 813
rect 2102 745 2136 779
rect 2068 711 2136 745
rect 2102 677 2136 711
rect 2068 643 2136 677
rect 2102 609 2136 643
rect 2068 575 2136 609
rect 2102 541 2136 575
rect 2068 507 2136 541
rect 2102 473 2136 507
rect 2068 439 2136 473
rect 2102 405 2136 439
rect 2068 371 2136 405
rect 2102 337 2136 371
rect 2068 303 2136 337
rect 2102 269 2136 303
rect 2068 235 2136 269
rect 2102 201 2136 235
rect 2238 201 2257 1595
rect 2068 185 2257 201
rect 190 163 230 185
rect 2068 163 2108 185
rect 190 147 256 163
rect 190 113 206 147
rect 240 113 256 147
rect 2042 147 2108 163
rect 190 97 256 113
rect 385 125 1913 137
rect 385 19 412 125
rect 1886 19 1913 125
rect 2042 113 2058 147
rect 2092 113 2108 147
rect 2042 97 2108 113
rect 385 0 1913 19
<< viali >>
rect 412 1775 1886 1777
rect 412 1673 418 1775
rect 418 1673 1880 1775
rect 1880 1673 1886 1775
rect 412 1671 1886 1673
rect 60 1529 94 1563
rect 60 1457 94 1491
rect 60 1385 94 1419
rect 60 1313 94 1347
rect 60 1241 94 1275
rect 60 1169 94 1203
rect 60 1097 94 1131
rect 60 1025 94 1059
rect 60 953 94 987
rect 60 881 94 915
rect 60 809 94 843
rect 60 737 94 771
rect 60 665 94 699
rect 60 593 94 627
rect 60 521 94 555
rect 60 449 94 483
rect 60 377 94 411
rect 60 305 94 339
rect 60 233 94 267
rect 352 1561 386 1563
rect 352 1529 386 1561
rect 352 1459 386 1491
rect 352 1457 386 1459
rect 352 1391 386 1419
rect 352 1385 386 1391
rect 352 1323 386 1347
rect 352 1313 386 1323
rect 352 1255 386 1275
rect 352 1241 386 1255
rect 352 1187 386 1203
rect 352 1169 386 1187
rect 352 1119 386 1131
rect 352 1097 386 1119
rect 352 1051 386 1059
rect 352 1025 386 1051
rect 352 983 386 987
rect 352 953 386 983
rect 352 881 386 915
rect 352 813 386 843
rect 352 809 386 813
rect 352 745 386 771
rect 352 737 386 745
rect 352 677 386 699
rect 352 665 386 677
rect 352 609 386 627
rect 352 593 386 609
rect 352 541 386 555
rect 352 521 386 541
rect 352 473 386 483
rect 352 449 386 473
rect 352 405 386 411
rect 352 377 386 405
rect 352 337 386 339
rect 352 305 386 337
rect 352 235 386 267
rect 352 233 386 235
rect 508 1561 542 1563
rect 508 1529 542 1561
rect 508 1459 542 1491
rect 508 1457 542 1459
rect 508 1391 542 1419
rect 508 1385 542 1391
rect 508 1323 542 1347
rect 508 1313 542 1323
rect 508 1255 542 1275
rect 508 1241 542 1255
rect 508 1187 542 1203
rect 508 1169 542 1187
rect 508 1119 542 1131
rect 508 1097 542 1119
rect 508 1051 542 1059
rect 508 1025 542 1051
rect 508 983 542 987
rect 508 953 542 983
rect 508 881 542 915
rect 508 813 542 843
rect 508 809 542 813
rect 508 745 542 771
rect 508 737 542 745
rect 508 677 542 699
rect 508 665 542 677
rect 508 609 542 627
rect 508 593 542 609
rect 508 541 542 555
rect 508 521 542 541
rect 508 473 542 483
rect 508 449 542 473
rect 508 405 542 411
rect 508 377 542 405
rect 508 337 542 339
rect 508 305 542 337
rect 508 235 542 267
rect 508 233 542 235
rect 664 1561 698 1563
rect 664 1529 698 1561
rect 664 1459 698 1491
rect 664 1457 698 1459
rect 664 1391 698 1419
rect 664 1385 698 1391
rect 664 1323 698 1347
rect 664 1313 698 1323
rect 664 1255 698 1275
rect 664 1241 698 1255
rect 664 1187 698 1203
rect 664 1169 698 1187
rect 664 1119 698 1131
rect 664 1097 698 1119
rect 664 1051 698 1059
rect 664 1025 698 1051
rect 664 983 698 987
rect 664 953 698 983
rect 664 881 698 915
rect 664 813 698 843
rect 664 809 698 813
rect 664 745 698 771
rect 664 737 698 745
rect 664 677 698 699
rect 664 665 698 677
rect 664 609 698 627
rect 664 593 698 609
rect 664 541 698 555
rect 664 521 698 541
rect 664 473 698 483
rect 664 449 698 473
rect 664 405 698 411
rect 664 377 698 405
rect 664 337 698 339
rect 664 305 698 337
rect 664 235 698 267
rect 664 233 698 235
rect 820 1561 854 1563
rect 820 1529 854 1561
rect 820 1459 854 1491
rect 820 1457 854 1459
rect 820 1391 854 1419
rect 820 1385 854 1391
rect 820 1323 854 1347
rect 820 1313 854 1323
rect 820 1255 854 1275
rect 820 1241 854 1255
rect 820 1187 854 1203
rect 820 1169 854 1187
rect 820 1119 854 1131
rect 820 1097 854 1119
rect 820 1051 854 1059
rect 820 1025 854 1051
rect 820 983 854 987
rect 820 953 854 983
rect 820 881 854 915
rect 820 813 854 843
rect 820 809 854 813
rect 820 745 854 771
rect 820 737 854 745
rect 820 677 854 699
rect 820 665 854 677
rect 820 609 854 627
rect 820 593 854 609
rect 820 541 854 555
rect 820 521 854 541
rect 820 473 854 483
rect 820 449 854 473
rect 820 405 854 411
rect 820 377 854 405
rect 820 337 854 339
rect 820 305 854 337
rect 820 235 854 267
rect 820 233 854 235
rect 976 1561 1010 1563
rect 976 1529 1010 1561
rect 976 1459 1010 1491
rect 976 1457 1010 1459
rect 976 1391 1010 1419
rect 976 1385 1010 1391
rect 976 1323 1010 1347
rect 976 1313 1010 1323
rect 976 1255 1010 1275
rect 976 1241 1010 1255
rect 976 1187 1010 1203
rect 976 1169 1010 1187
rect 976 1119 1010 1131
rect 976 1097 1010 1119
rect 976 1051 1010 1059
rect 976 1025 1010 1051
rect 976 983 1010 987
rect 976 953 1010 983
rect 976 881 1010 915
rect 976 813 1010 843
rect 976 809 1010 813
rect 976 745 1010 771
rect 976 737 1010 745
rect 976 677 1010 699
rect 976 665 1010 677
rect 976 609 1010 627
rect 976 593 1010 609
rect 976 541 1010 555
rect 976 521 1010 541
rect 976 473 1010 483
rect 976 449 1010 473
rect 976 405 1010 411
rect 976 377 1010 405
rect 976 337 1010 339
rect 976 305 1010 337
rect 976 235 1010 267
rect 976 233 1010 235
rect 1132 1561 1166 1563
rect 1132 1529 1166 1561
rect 1132 1459 1166 1491
rect 1132 1457 1166 1459
rect 1132 1391 1166 1419
rect 1132 1385 1166 1391
rect 1132 1323 1166 1347
rect 1132 1313 1166 1323
rect 1132 1255 1166 1275
rect 1132 1241 1166 1255
rect 1132 1187 1166 1203
rect 1132 1169 1166 1187
rect 1132 1119 1166 1131
rect 1132 1097 1166 1119
rect 1132 1051 1166 1059
rect 1132 1025 1166 1051
rect 1132 983 1166 987
rect 1132 953 1166 983
rect 1132 881 1166 915
rect 1132 813 1166 843
rect 1132 809 1166 813
rect 1132 745 1166 771
rect 1132 737 1166 745
rect 1132 677 1166 699
rect 1132 665 1166 677
rect 1132 609 1166 627
rect 1132 593 1166 609
rect 1132 541 1166 555
rect 1132 521 1166 541
rect 1132 473 1166 483
rect 1132 449 1166 473
rect 1132 405 1166 411
rect 1132 377 1166 405
rect 1132 337 1166 339
rect 1132 305 1166 337
rect 1132 235 1166 267
rect 1132 233 1166 235
rect 1288 1561 1322 1563
rect 1288 1529 1322 1561
rect 1288 1459 1322 1491
rect 1288 1457 1322 1459
rect 1288 1391 1322 1419
rect 1288 1385 1322 1391
rect 1288 1323 1322 1347
rect 1288 1313 1322 1323
rect 1288 1255 1322 1275
rect 1288 1241 1322 1255
rect 1288 1187 1322 1203
rect 1288 1169 1322 1187
rect 1288 1119 1322 1131
rect 1288 1097 1322 1119
rect 1288 1051 1322 1059
rect 1288 1025 1322 1051
rect 1288 983 1322 987
rect 1288 953 1322 983
rect 1288 881 1322 915
rect 1288 813 1322 843
rect 1288 809 1322 813
rect 1288 745 1322 771
rect 1288 737 1322 745
rect 1288 677 1322 699
rect 1288 665 1322 677
rect 1288 609 1322 627
rect 1288 593 1322 609
rect 1288 541 1322 555
rect 1288 521 1322 541
rect 1288 473 1322 483
rect 1288 449 1322 473
rect 1288 405 1322 411
rect 1288 377 1322 405
rect 1288 337 1322 339
rect 1288 305 1322 337
rect 1288 235 1322 267
rect 1288 233 1322 235
rect 1444 1561 1478 1563
rect 1444 1529 1478 1561
rect 1444 1459 1478 1491
rect 1444 1457 1478 1459
rect 1444 1391 1478 1419
rect 1444 1385 1478 1391
rect 1444 1323 1478 1347
rect 1444 1313 1478 1323
rect 1444 1255 1478 1275
rect 1444 1241 1478 1255
rect 1444 1187 1478 1203
rect 1444 1169 1478 1187
rect 1444 1119 1478 1131
rect 1444 1097 1478 1119
rect 1444 1051 1478 1059
rect 1444 1025 1478 1051
rect 1444 983 1478 987
rect 1444 953 1478 983
rect 1444 881 1478 915
rect 1444 813 1478 843
rect 1444 809 1478 813
rect 1444 745 1478 771
rect 1444 737 1478 745
rect 1444 677 1478 699
rect 1444 665 1478 677
rect 1444 609 1478 627
rect 1444 593 1478 609
rect 1444 541 1478 555
rect 1444 521 1478 541
rect 1444 473 1478 483
rect 1444 449 1478 473
rect 1444 405 1478 411
rect 1444 377 1478 405
rect 1444 337 1478 339
rect 1444 305 1478 337
rect 1444 235 1478 267
rect 1444 233 1478 235
rect 1600 1561 1634 1563
rect 1600 1529 1634 1561
rect 1600 1459 1634 1491
rect 1600 1457 1634 1459
rect 1600 1391 1634 1419
rect 1600 1385 1634 1391
rect 1600 1323 1634 1347
rect 1600 1313 1634 1323
rect 1600 1255 1634 1275
rect 1600 1241 1634 1255
rect 1600 1187 1634 1203
rect 1600 1169 1634 1187
rect 1600 1119 1634 1131
rect 1600 1097 1634 1119
rect 1600 1051 1634 1059
rect 1600 1025 1634 1051
rect 1600 983 1634 987
rect 1600 953 1634 983
rect 1600 881 1634 915
rect 1600 813 1634 843
rect 1600 809 1634 813
rect 1600 745 1634 771
rect 1600 737 1634 745
rect 1600 677 1634 699
rect 1600 665 1634 677
rect 1600 609 1634 627
rect 1600 593 1634 609
rect 1600 541 1634 555
rect 1600 521 1634 541
rect 1600 473 1634 483
rect 1600 449 1634 473
rect 1600 405 1634 411
rect 1600 377 1634 405
rect 1600 337 1634 339
rect 1600 305 1634 337
rect 1600 235 1634 267
rect 1600 233 1634 235
rect 1756 1561 1790 1563
rect 1756 1529 1790 1561
rect 1756 1459 1790 1491
rect 1756 1457 1790 1459
rect 1756 1391 1790 1419
rect 1756 1385 1790 1391
rect 1756 1323 1790 1347
rect 1756 1313 1790 1323
rect 1756 1255 1790 1275
rect 1756 1241 1790 1255
rect 1756 1187 1790 1203
rect 1756 1169 1790 1187
rect 1756 1119 1790 1131
rect 1756 1097 1790 1119
rect 1756 1051 1790 1059
rect 1756 1025 1790 1051
rect 1756 983 1790 987
rect 1756 953 1790 983
rect 1756 881 1790 915
rect 1756 813 1790 843
rect 1756 809 1790 813
rect 1756 745 1790 771
rect 1756 737 1790 745
rect 1756 677 1790 699
rect 1756 665 1790 677
rect 1756 609 1790 627
rect 1756 593 1790 609
rect 1756 541 1790 555
rect 1756 521 1790 541
rect 1756 473 1790 483
rect 1756 449 1790 473
rect 1756 405 1790 411
rect 1756 377 1790 405
rect 1756 337 1790 339
rect 1756 305 1790 337
rect 1756 235 1790 267
rect 1756 233 1790 235
rect 1912 1561 1946 1563
rect 1912 1529 1946 1561
rect 1912 1459 1946 1491
rect 1912 1457 1946 1459
rect 1912 1391 1946 1419
rect 1912 1385 1946 1391
rect 1912 1323 1946 1347
rect 1912 1313 1946 1323
rect 1912 1255 1946 1275
rect 1912 1241 1946 1255
rect 1912 1187 1946 1203
rect 1912 1169 1946 1187
rect 1912 1119 1946 1131
rect 1912 1097 1946 1119
rect 1912 1051 1946 1059
rect 1912 1025 1946 1051
rect 1912 983 1946 987
rect 1912 953 1946 983
rect 1912 881 1946 915
rect 1912 813 1946 843
rect 1912 809 1946 813
rect 1912 745 1946 771
rect 1912 737 1946 745
rect 1912 677 1946 699
rect 1912 665 1946 677
rect 1912 609 1946 627
rect 1912 593 1946 609
rect 1912 541 1946 555
rect 1912 521 1946 541
rect 1912 473 1946 483
rect 1912 449 1946 473
rect 1912 405 1946 411
rect 1912 377 1946 405
rect 1912 337 1946 339
rect 1912 305 1946 337
rect 1912 235 1946 267
rect 1912 233 1946 235
rect 2204 1529 2238 1563
rect 2204 1457 2238 1491
rect 2204 1385 2238 1419
rect 2204 1313 2238 1347
rect 2204 1241 2238 1275
rect 2204 1169 2238 1203
rect 2204 1097 2238 1131
rect 2204 1025 2238 1059
rect 2204 953 2238 987
rect 2204 881 2238 915
rect 2204 809 2238 843
rect 2204 737 2238 771
rect 2204 665 2238 699
rect 2204 593 2238 627
rect 2204 521 2238 555
rect 2204 449 2238 483
rect 2204 377 2238 411
rect 2204 305 2238 339
rect 2204 233 2238 267
rect 412 123 1886 125
rect 412 21 418 123
rect 418 21 1880 123
rect 1880 21 1886 123
rect 412 19 1886 21
<< metal1 >>
rect 381 1777 1917 1796
rect 381 1671 412 1777
rect 1886 1671 1917 1777
rect 381 1659 1917 1671
rect 41 1563 100 1594
rect 41 1529 60 1563
rect 94 1529 100 1563
rect 41 1491 100 1529
rect 41 1457 60 1491
rect 94 1457 100 1491
rect 41 1419 100 1457
rect 41 1385 60 1419
rect 94 1385 100 1419
rect 41 1347 100 1385
rect 41 1313 60 1347
rect 94 1313 100 1347
rect 41 1275 100 1313
rect 41 1241 60 1275
rect 94 1241 100 1275
rect 41 1203 100 1241
rect 41 1169 60 1203
rect 94 1169 100 1203
rect 41 1131 100 1169
rect 41 1097 60 1131
rect 94 1097 100 1131
rect 41 1059 100 1097
rect 41 1025 60 1059
rect 94 1025 100 1059
rect 41 987 100 1025
rect 41 953 60 987
rect 94 953 100 987
rect 41 915 100 953
rect 41 881 60 915
rect 94 881 100 915
rect 41 843 100 881
rect 41 809 60 843
rect 94 809 100 843
rect 41 771 100 809
rect 41 737 60 771
rect 94 737 100 771
rect 41 699 100 737
rect 41 665 60 699
rect 94 665 100 699
rect 41 627 100 665
rect 41 593 60 627
rect 94 593 100 627
rect 41 555 100 593
rect 41 521 60 555
rect 94 521 100 555
rect 41 483 100 521
rect 41 449 60 483
rect 94 449 100 483
rect 41 411 100 449
rect 41 377 60 411
rect 94 377 100 411
rect 41 339 100 377
rect 41 305 60 339
rect 94 305 100 339
rect 41 267 100 305
rect 41 233 60 267
rect 94 233 100 267
rect 41 202 100 233
rect 343 1588 395 1594
rect 343 1529 352 1536
rect 386 1529 395 1536
rect 343 1524 395 1529
rect 343 1460 352 1472
rect 386 1460 395 1472
rect 343 1396 352 1408
rect 386 1396 395 1408
rect 343 1332 352 1344
rect 386 1332 395 1344
rect 343 1275 395 1280
rect 343 1241 352 1275
rect 386 1241 395 1275
rect 343 1203 395 1241
rect 343 1169 352 1203
rect 386 1169 395 1203
rect 343 1131 395 1169
rect 343 1097 352 1131
rect 386 1097 395 1131
rect 343 1059 395 1097
rect 343 1025 352 1059
rect 386 1025 395 1059
rect 343 987 395 1025
rect 343 953 352 987
rect 386 953 395 987
rect 343 915 395 953
rect 343 881 352 915
rect 386 881 395 915
rect 343 843 395 881
rect 343 809 352 843
rect 386 809 395 843
rect 343 771 395 809
rect 343 737 352 771
rect 386 737 395 771
rect 343 699 395 737
rect 343 665 352 699
rect 386 665 395 699
rect 343 627 395 665
rect 343 593 352 627
rect 386 593 395 627
rect 343 555 395 593
rect 343 521 352 555
rect 386 521 395 555
rect 343 516 395 521
rect 343 452 352 464
rect 386 452 395 464
rect 343 388 352 400
rect 386 388 395 400
rect 343 324 352 336
rect 386 324 395 336
rect 343 267 395 272
rect 343 260 352 267
rect 386 260 395 267
rect 343 202 395 208
rect 499 1563 551 1594
rect 499 1529 508 1563
rect 542 1529 551 1563
rect 499 1491 551 1529
rect 499 1457 508 1491
rect 542 1457 551 1491
rect 499 1419 551 1457
rect 499 1385 508 1419
rect 542 1385 551 1419
rect 499 1347 551 1385
rect 499 1313 508 1347
rect 542 1313 551 1347
rect 499 1275 551 1313
rect 499 1241 508 1275
rect 542 1241 551 1275
rect 499 1212 551 1241
rect 499 1148 551 1160
rect 499 1084 551 1096
rect 499 1025 508 1032
rect 542 1025 551 1032
rect 499 1020 551 1025
rect 499 956 508 968
rect 542 956 551 968
rect 499 892 508 904
rect 542 892 551 904
rect 499 828 508 840
rect 542 828 551 840
rect 499 771 551 776
rect 499 764 508 771
rect 542 764 551 771
rect 499 700 551 712
rect 499 636 551 648
rect 499 555 551 584
rect 499 521 508 555
rect 542 521 551 555
rect 499 483 551 521
rect 499 449 508 483
rect 542 449 551 483
rect 499 411 551 449
rect 499 377 508 411
rect 542 377 551 411
rect 499 339 551 377
rect 499 305 508 339
rect 542 305 551 339
rect 499 267 551 305
rect 499 233 508 267
rect 542 233 551 267
rect 499 202 551 233
rect 655 1588 707 1594
rect 655 1529 664 1536
rect 698 1529 707 1536
rect 655 1524 707 1529
rect 655 1460 664 1472
rect 698 1460 707 1472
rect 655 1396 664 1408
rect 698 1396 707 1408
rect 655 1332 664 1344
rect 698 1332 707 1344
rect 655 1275 707 1280
rect 655 1241 664 1275
rect 698 1241 707 1275
rect 655 1203 707 1241
rect 655 1169 664 1203
rect 698 1169 707 1203
rect 655 1131 707 1169
rect 655 1097 664 1131
rect 698 1097 707 1131
rect 655 1059 707 1097
rect 655 1025 664 1059
rect 698 1025 707 1059
rect 655 987 707 1025
rect 655 953 664 987
rect 698 953 707 987
rect 655 915 707 953
rect 655 881 664 915
rect 698 881 707 915
rect 655 843 707 881
rect 655 809 664 843
rect 698 809 707 843
rect 655 771 707 809
rect 655 737 664 771
rect 698 737 707 771
rect 655 699 707 737
rect 655 665 664 699
rect 698 665 707 699
rect 655 627 707 665
rect 655 593 664 627
rect 698 593 707 627
rect 655 555 707 593
rect 655 521 664 555
rect 698 521 707 555
rect 655 516 707 521
rect 655 452 664 464
rect 698 452 707 464
rect 655 388 664 400
rect 698 388 707 400
rect 655 324 664 336
rect 698 324 707 336
rect 655 267 707 272
rect 655 260 664 267
rect 698 260 707 267
rect 655 202 707 208
rect 811 1563 863 1594
rect 811 1529 820 1563
rect 854 1529 863 1563
rect 811 1491 863 1529
rect 811 1457 820 1491
rect 854 1457 863 1491
rect 811 1419 863 1457
rect 811 1385 820 1419
rect 854 1385 863 1419
rect 811 1347 863 1385
rect 811 1313 820 1347
rect 854 1313 863 1347
rect 811 1275 863 1313
rect 811 1241 820 1275
rect 854 1241 863 1275
rect 811 1212 863 1241
rect 811 1148 863 1160
rect 811 1084 863 1096
rect 811 1025 820 1032
rect 854 1025 863 1032
rect 811 1020 863 1025
rect 811 956 820 968
rect 854 956 863 968
rect 811 892 820 904
rect 854 892 863 904
rect 811 828 820 840
rect 854 828 863 840
rect 811 771 863 776
rect 811 764 820 771
rect 854 764 863 771
rect 811 700 863 712
rect 811 636 863 648
rect 811 555 863 584
rect 811 521 820 555
rect 854 521 863 555
rect 811 483 863 521
rect 811 449 820 483
rect 854 449 863 483
rect 811 411 863 449
rect 811 377 820 411
rect 854 377 863 411
rect 811 339 863 377
rect 811 305 820 339
rect 854 305 863 339
rect 811 267 863 305
rect 811 233 820 267
rect 854 233 863 267
rect 811 202 863 233
rect 967 1588 1019 1594
rect 967 1529 976 1536
rect 1010 1529 1019 1536
rect 967 1524 1019 1529
rect 967 1460 976 1472
rect 1010 1460 1019 1472
rect 967 1396 976 1408
rect 1010 1396 1019 1408
rect 967 1332 976 1344
rect 1010 1332 1019 1344
rect 967 1275 1019 1280
rect 967 1241 976 1275
rect 1010 1241 1019 1275
rect 967 1203 1019 1241
rect 967 1169 976 1203
rect 1010 1169 1019 1203
rect 967 1131 1019 1169
rect 967 1097 976 1131
rect 1010 1097 1019 1131
rect 967 1059 1019 1097
rect 967 1025 976 1059
rect 1010 1025 1019 1059
rect 967 987 1019 1025
rect 967 953 976 987
rect 1010 953 1019 987
rect 967 915 1019 953
rect 967 881 976 915
rect 1010 881 1019 915
rect 967 843 1019 881
rect 967 809 976 843
rect 1010 809 1019 843
rect 967 771 1019 809
rect 967 737 976 771
rect 1010 737 1019 771
rect 967 699 1019 737
rect 967 665 976 699
rect 1010 665 1019 699
rect 967 627 1019 665
rect 967 593 976 627
rect 1010 593 1019 627
rect 967 555 1019 593
rect 967 521 976 555
rect 1010 521 1019 555
rect 967 516 1019 521
rect 967 452 976 464
rect 1010 452 1019 464
rect 967 388 976 400
rect 1010 388 1019 400
rect 967 324 976 336
rect 1010 324 1019 336
rect 967 267 1019 272
rect 967 260 976 267
rect 1010 260 1019 267
rect 967 202 1019 208
rect 1123 1563 1175 1594
rect 1123 1529 1132 1563
rect 1166 1529 1175 1563
rect 1123 1491 1175 1529
rect 1123 1457 1132 1491
rect 1166 1457 1175 1491
rect 1123 1419 1175 1457
rect 1123 1385 1132 1419
rect 1166 1385 1175 1419
rect 1123 1347 1175 1385
rect 1123 1313 1132 1347
rect 1166 1313 1175 1347
rect 1123 1275 1175 1313
rect 1123 1241 1132 1275
rect 1166 1241 1175 1275
rect 1123 1212 1175 1241
rect 1123 1148 1175 1160
rect 1123 1084 1175 1096
rect 1123 1025 1132 1032
rect 1166 1025 1175 1032
rect 1123 1020 1175 1025
rect 1123 956 1132 968
rect 1166 956 1175 968
rect 1123 892 1132 904
rect 1166 892 1175 904
rect 1123 828 1132 840
rect 1166 828 1175 840
rect 1123 771 1175 776
rect 1123 764 1132 771
rect 1166 764 1175 771
rect 1123 700 1175 712
rect 1123 636 1175 648
rect 1123 555 1175 584
rect 1123 521 1132 555
rect 1166 521 1175 555
rect 1123 483 1175 521
rect 1123 449 1132 483
rect 1166 449 1175 483
rect 1123 411 1175 449
rect 1123 377 1132 411
rect 1166 377 1175 411
rect 1123 339 1175 377
rect 1123 305 1132 339
rect 1166 305 1175 339
rect 1123 267 1175 305
rect 1123 233 1132 267
rect 1166 233 1175 267
rect 1123 202 1175 233
rect 1279 1588 1331 1594
rect 1279 1529 1288 1536
rect 1322 1529 1331 1536
rect 1279 1524 1331 1529
rect 1279 1460 1288 1472
rect 1322 1460 1331 1472
rect 1279 1396 1288 1408
rect 1322 1396 1331 1408
rect 1279 1332 1288 1344
rect 1322 1332 1331 1344
rect 1279 1275 1331 1280
rect 1279 1241 1288 1275
rect 1322 1241 1331 1275
rect 1279 1203 1331 1241
rect 1279 1169 1288 1203
rect 1322 1169 1331 1203
rect 1279 1131 1331 1169
rect 1279 1097 1288 1131
rect 1322 1097 1331 1131
rect 1279 1059 1331 1097
rect 1279 1025 1288 1059
rect 1322 1025 1331 1059
rect 1279 987 1331 1025
rect 1279 953 1288 987
rect 1322 953 1331 987
rect 1279 915 1331 953
rect 1279 881 1288 915
rect 1322 881 1331 915
rect 1279 843 1331 881
rect 1279 809 1288 843
rect 1322 809 1331 843
rect 1279 771 1331 809
rect 1279 737 1288 771
rect 1322 737 1331 771
rect 1279 699 1331 737
rect 1279 665 1288 699
rect 1322 665 1331 699
rect 1279 627 1331 665
rect 1279 593 1288 627
rect 1322 593 1331 627
rect 1279 555 1331 593
rect 1279 521 1288 555
rect 1322 521 1331 555
rect 1279 516 1331 521
rect 1279 452 1288 464
rect 1322 452 1331 464
rect 1279 388 1288 400
rect 1322 388 1331 400
rect 1279 324 1288 336
rect 1322 324 1331 336
rect 1279 267 1331 272
rect 1279 260 1288 267
rect 1322 260 1331 267
rect 1279 202 1331 208
rect 1435 1563 1487 1594
rect 1435 1529 1444 1563
rect 1478 1529 1487 1563
rect 1435 1491 1487 1529
rect 1435 1457 1444 1491
rect 1478 1457 1487 1491
rect 1435 1419 1487 1457
rect 1435 1385 1444 1419
rect 1478 1385 1487 1419
rect 1435 1347 1487 1385
rect 1435 1313 1444 1347
rect 1478 1313 1487 1347
rect 1435 1275 1487 1313
rect 1435 1241 1444 1275
rect 1478 1241 1487 1275
rect 1435 1212 1487 1241
rect 1435 1148 1487 1160
rect 1435 1084 1487 1096
rect 1435 1025 1444 1032
rect 1478 1025 1487 1032
rect 1435 1020 1487 1025
rect 1435 956 1444 968
rect 1478 956 1487 968
rect 1435 892 1444 904
rect 1478 892 1487 904
rect 1435 828 1444 840
rect 1478 828 1487 840
rect 1435 771 1487 776
rect 1435 764 1444 771
rect 1478 764 1487 771
rect 1435 700 1487 712
rect 1435 636 1487 648
rect 1435 555 1487 584
rect 1435 521 1444 555
rect 1478 521 1487 555
rect 1435 483 1487 521
rect 1435 449 1444 483
rect 1478 449 1487 483
rect 1435 411 1487 449
rect 1435 377 1444 411
rect 1478 377 1487 411
rect 1435 339 1487 377
rect 1435 305 1444 339
rect 1478 305 1487 339
rect 1435 267 1487 305
rect 1435 233 1444 267
rect 1478 233 1487 267
rect 1435 202 1487 233
rect 1591 1588 1643 1594
rect 1591 1529 1600 1536
rect 1634 1529 1643 1536
rect 1591 1524 1643 1529
rect 1591 1460 1600 1472
rect 1634 1460 1643 1472
rect 1591 1396 1600 1408
rect 1634 1396 1643 1408
rect 1591 1332 1600 1344
rect 1634 1332 1643 1344
rect 1591 1275 1643 1280
rect 1591 1241 1600 1275
rect 1634 1241 1643 1275
rect 1591 1203 1643 1241
rect 1591 1169 1600 1203
rect 1634 1169 1643 1203
rect 1591 1131 1643 1169
rect 1591 1097 1600 1131
rect 1634 1097 1643 1131
rect 1591 1059 1643 1097
rect 1591 1025 1600 1059
rect 1634 1025 1643 1059
rect 1591 987 1643 1025
rect 1591 953 1600 987
rect 1634 953 1643 987
rect 1591 915 1643 953
rect 1591 881 1600 915
rect 1634 881 1643 915
rect 1591 843 1643 881
rect 1591 809 1600 843
rect 1634 809 1643 843
rect 1591 771 1643 809
rect 1591 737 1600 771
rect 1634 737 1643 771
rect 1591 699 1643 737
rect 1591 665 1600 699
rect 1634 665 1643 699
rect 1591 627 1643 665
rect 1591 593 1600 627
rect 1634 593 1643 627
rect 1591 555 1643 593
rect 1591 521 1600 555
rect 1634 521 1643 555
rect 1591 516 1643 521
rect 1591 452 1600 464
rect 1634 452 1643 464
rect 1591 388 1600 400
rect 1634 388 1643 400
rect 1591 324 1600 336
rect 1634 324 1643 336
rect 1591 267 1643 272
rect 1591 260 1600 267
rect 1634 260 1643 267
rect 1591 202 1643 208
rect 1747 1563 1799 1594
rect 1747 1529 1756 1563
rect 1790 1529 1799 1563
rect 1747 1491 1799 1529
rect 1747 1457 1756 1491
rect 1790 1457 1799 1491
rect 1747 1419 1799 1457
rect 1747 1385 1756 1419
rect 1790 1385 1799 1419
rect 1747 1347 1799 1385
rect 1747 1313 1756 1347
rect 1790 1313 1799 1347
rect 1747 1275 1799 1313
rect 1747 1241 1756 1275
rect 1790 1241 1799 1275
rect 1747 1212 1799 1241
rect 1747 1148 1799 1160
rect 1747 1084 1799 1096
rect 1747 1025 1756 1032
rect 1790 1025 1799 1032
rect 1747 1020 1799 1025
rect 1747 956 1756 968
rect 1790 956 1799 968
rect 1747 892 1756 904
rect 1790 892 1799 904
rect 1747 828 1756 840
rect 1790 828 1799 840
rect 1747 771 1799 776
rect 1747 764 1756 771
rect 1790 764 1799 771
rect 1747 700 1799 712
rect 1747 636 1799 648
rect 1747 555 1799 584
rect 1747 521 1756 555
rect 1790 521 1799 555
rect 1747 483 1799 521
rect 1747 449 1756 483
rect 1790 449 1799 483
rect 1747 411 1799 449
rect 1747 377 1756 411
rect 1790 377 1799 411
rect 1747 339 1799 377
rect 1747 305 1756 339
rect 1790 305 1799 339
rect 1747 267 1799 305
rect 1747 233 1756 267
rect 1790 233 1799 267
rect 1747 202 1799 233
rect 1903 1588 1955 1594
rect 1903 1529 1912 1536
rect 1946 1529 1955 1536
rect 1903 1524 1955 1529
rect 1903 1460 1912 1472
rect 1946 1460 1955 1472
rect 1903 1396 1912 1408
rect 1946 1396 1955 1408
rect 1903 1332 1912 1344
rect 1946 1332 1955 1344
rect 1903 1275 1955 1280
rect 1903 1241 1912 1275
rect 1946 1241 1955 1275
rect 1903 1203 1955 1241
rect 1903 1169 1912 1203
rect 1946 1169 1955 1203
rect 1903 1131 1955 1169
rect 1903 1097 1912 1131
rect 1946 1097 1955 1131
rect 1903 1059 1955 1097
rect 1903 1025 1912 1059
rect 1946 1025 1955 1059
rect 1903 987 1955 1025
rect 1903 953 1912 987
rect 1946 953 1955 987
rect 1903 915 1955 953
rect 1903 881 1912 915
rect 1946 881 1955 915
rect 1903 843 1955 881
rect 1903 809 1912 843
rect 1946 809 1955 843
rect 1903 771 1955 809
rect 1903 737 1912 771
rect 1946 737 1955 771
rect 1903 699 1955 737
rect 1903 665 1912 699
rect 1946 665 1955 699
rect 1903 627 1955 665
rect 1903 593 1912 627
rect 1946 593 1955 627
rect 1903 555 1955 593
rect 1903 521 1912 555
rect 1946 521 1955 555
rect 1903 516 1955 521
rect 1903 452 1912 464
rect 1946 452 1955 464
rect 1903 388 1912 400
rect 1946 388 1955 400
rect 1903 324 1912 336
rect 1946 324 1955 336
rect 1903 267 1955 272
rect 1903 260 1912 267
rect 1946 260 1955 267
rect 1903 202 1955 208
rect 2198 1563 2257 1594
rect 2198 1529 2204 1563
rect 2238 1529 2257 1563
rect 2198 1491 2257 1529
rect 2198 1457 2204 1491
rect 2238 1457 2257 1491
rect 2198 1419 2257 1457
rect 2198 1385 2204 1419
rect 2238 1385 2257 1419
rect 2198 1347 2257 1385
rect 2198 1313 2204 1347
rect 2238 1313 2257 1347
rect 2198 1275 2257 1313
rect 2198 1241 2204 1275
rect 2238 1241 2257 1275
rect 2198 1203 2257 1241
rect 2198 1169 2204 1203
rect 2238 1169 2257 1203
rect 2198 1131 2257 1169
rect 2198 1097 2204 1131
rect 2238 1097 2257 1131
rect 2198 1059 2257 1097
rect 2198 1025 2204 1059
rect 2238 1025 2257 1059
rect 2198 987 2257 1025
rect 2198 953 2204 987
rect 2238 953 2257 987
rect 2198 915 2257 953
rect 2198 881 2204 915
rect 2238 881 2257 915
rect 2198 843 2257 881
rect 2198 809 2204 843
rect 2238 809 2257 843
rect 2198 771 2257 809
rect 2198 737 2204 771
rect 2238 737 2257 771
rect 2198 699 2257 737
rect 2198 665 2204 699
rect 2238 665 2257 699
rect 2198 627 2257 665
rect 2198 593 2204 627
rect 2238 593 2257 627
rect 2198 555 2257 593
rect 2198 521 2204 555
rect 2238 521 2257 555
rect 2198 483 2257 521
rect 2198 449 2204 483
rect 2238 449 2257 483
rect 2198 411 2257 449
rect 2198 377 2204 411
rect 2238 377 2257 411
rect 2198 339 2257 377
rect 2198 305 2204 339
rect 2238 305 2257 339
rect 2198 267 2257 305
rect 2198 233 2204 267
rect 2238 233 2257 267
rect 2198 202 2257 233
rect 381 125 1917 137
rect 381 19 412 125
rect 1886 19 1917 125
rect 381 0 1917 19
<< via1 >>
rect 343 1563 395 1588
rect 343 1536 352 1563
rect 352 1536 386 1563
rect 386 1536 395 1563
rect 343 1491 395 1524
rect 343 1472 352 1491
rect 352 1472 386 1491
rect 386 1472 395 1491
rect 343 1457 352 1460
rect 352 1457 386 1460
rect 386 1457 395 1460
rect 343 1419 395 1457
rect 343 1408 352 1419
rect 352 1408 386 1419
rect 386 1408 395 1419
rect 343 1385 352 1396
rect 352 1385 386 1396
rect 386 1385 395 1396
rect 343 1347 395 1385
rect 343 1344 352 1347
rect 352 1344 386 1347
rect 386 1344 395 1347
rect 343 1313 352 1332
rect 352 1313 386 1332
rect 386 1313 395 1332
rect 343 1280 395 1313
rect 343 483 395 516
rect 343 464 352 483
rect 352 464 386 483
rect 386 464 395 483
rect 343 449 352 452
rect 352 449 386 452
rect 386 449 395 452
rect 343 411 395 449
rect 343 400 352 411
rect 352 400 386 411
rect 386 400 395 411
rect 343 377 352 388
rect 352 377 386 388
rect 386 377 395 388
rect 343 339 395 377
rect 343 336 352 339
rect 352 336 386 339
rect 386 336 395 339
rect 343 305 352 324
rect 352 305 386 324
rect 386 305 395 324
rect 343 272 395 305
rect 343 233 352 260
rect 352 233 386 260
rect 386 233 395 260
rect 343 208 395 233
rect 499 1203 551 1212
rect 499 1169 508 1203
rect 508 1169 542 1203
rect 542 1169 551 1203
rect 499 1160 551 1169
rect 499 1131 551 1148
rect 499 1097 508 1131
rect 508 1097 542 1131
rect 542 1097 551 1131
rect 499 1096 551 1097
rect 499 1059 551 1084
rect 499 1032 508 1059
rect 508 1032 542 1059
rect 542 1032 551 1059
rect 499 987 551 1020
rect 499 968 508 987
rect 508 968 542 987
rect 542 968 551 987
rect 499 953 508 956
rect 508 953 542 956
rect 542 953 551 956
rect 499 915 551 953
rect 499 904 508 915
rect 508 904 542 915
rect 542 904 551 915
rect 499 881 508 892
rect 508 881 542 892
rect 542 881 551 892
rect 499 843 551 881
rect 499 840 508 843
rect 508 840 542 843
rect 542 840 551 843
rect 499 809 508 828
rect 508 809 542 828
rect 542 809 551 828
rect 499 776 551 809
rect 499 737 508 764
rect 508 737 542 764
rect 542 737 551 764
rect 499 712 551 737
rect 499 699 551 700
rect 499 665 508 699
rect 508 665 542 699
rect 542 665 551 699
rect 499 648 551 665
rect 499 627 551 636
rect 499 593 508 627
rect 508 593 542 627
rect 542 593 551 627
rect 499 584 551 593
rect 655 1563 707 1588
rect 655 1536 664 1563
rect 664 1536 698 1563
rect 698 1536 707 1563
rect 655 1491 707 1524
rect 655 1472 664 1491
rect 664 1472 698 1491
rect 698 1472 707 1491
rect 655 1457 664 1460
rect 664 1457 698 1460
rect 698 1457 707 1460
rect 655 1419 707 1457
rect 655 1408 664 1419
rect 664 1408 698 1419
rect 698 1408 707 1419
rect 655 1385 664 1396
rect 664 1385 698 1396
rect 698 1385 707 1396
rect 655 1347 707 1385
rect 655 1344 664 1347
rect 664 1344 698 1347
rect 698 1344 707 1347
rect 655 1313 664 1332
rect 664 1313 698 1332
rect 698 1313 707 1332
rect 655 1280 707 1313
rect 655 483 707 516
rect 655 464 664 483
rect 664 464 698 483
rect 698 464 707 483
rect 655 449 664 452
rect 664 449 698 452
rect 698 449 707 452
rect 655 411 707 449
rect 655 400 664 411
rect 664 400 698 411
rect 698 400 707 411
rect 655 377 664 388
rect 664 377 698 388
rect 698 377 707 388
rect 655 339 707 377
rect 655 336 664 339
rect 664 336 698 339
rect 698 336 707 339
rect 655 305 664 324
rect 664 305 698 324
rect 698 305 707 324
rect 655 272 707 305
rect 655 233 664 260
rect 664 233 698 260
rect 698 233 707 260
rect 655 208 707 233
rect 811 1203 863 1212
rect 811 1169 820 1203
rect 820 1169 854 1203
rect 854 1169 863 1203
rect 811 1160 863 1169
rect 811 1131 863 1148
rect 811 1097 820 1131
rect 820 1097 854 1131
rect 854 1097 863 1131
rect 811 1096 863 1097
rect 811 1059 863 1084
rect 811 1032 820 1059
rect 820 1032 854 1059
rect 854 1032 863 1059
rect 811 987 863 1020
rect 811 968 820 987
rect 820 968 854 987
rect 854 968 863 987
rect 811 953 820 956
rect 820 953 854 956
rect 854 953 863 956
rect 811 915 863 953
rect 811 904 820 915
rect 820 904 854 915
rect 854 904 863 915
rect 811 881 820 892
rect 820 881 854 892
rect 854 881 863 892
rect 811 843 863 881
rect 811 840 820 843
rect 820 840 854 843
rect 854 840 863 843
rect 811 809 820 828
rect 820 809 854 828
rect 854 809 863 828
rect 811 776 863 809
rect 811 737 820 764
rect 820 737 854 764
rect 854 737 863 764
rect 811 712 863 737
rect 811 699 863 700
rect 811 665 820 699
rect 820 665 854 699
rect 854 665 863 699
rect 811 648 863 665
rect 811 627 863 636
rect 811 593 820 627
rect 820 593 854 627
rect 854 593 863 627
rect 811 584 863 593
rect 967 1563 1019 1588
rect 967 1536 976 1563
rect 976 1536 1010 1563
rect 1010 1536 1019 1563
rect 967 1491 1019 1524
rect 967 1472 976 1491
rect 976 1472 1010 1491
rect 1010 1472 1019 1491
rect 967 1457 976 1460
rect 976 1457 1010 1460
rect 1010 1457 1019 1460
rect 967 1419 1019 1457
rect 967 1408 976 1419
rect 976 1408 1010 1419
rect 1010 1408 1019 1419
rect 967 1385 976 1396
rect 976 1385 1010 1396
rect 1010 1385 1019 1396
rect 967 1347 1019 1385
rect 967 1344 976 1347
rect 976 1344 1010 1347
rect 1010 1344 1019 1347
rect 967 1313 976 1332
rect 976 1313 1010 1332
rect 1010 1313 1019 1332
rect 967 1280 1019 1313
rect 967 483 1019 516
rect 967 464 976 483
rect 976 464 1010 483
rect 1010 464 1019 483
rect 967 449 976 452
rect 976 449 1010 452
rect 1010 449 1019 452
rect 967 411 1019 449
rect 967 400 976 411
rect 976 400 1010 411
rect 1010 400 1019 411
rect 967 377 976 388
rect 976 377 1010 388
rect 1010 377 1019 388
rect 967 339 1019 377
rect 967 336 976 339
rect 976 336 1010 339
rect 1010 336 1019 339
rect 967 305 976 324
rect 976 305 1010 324
rect 1010 305 1019 324
rect 967 272 1019 305
rect 967 233 976 260
rect 976 233 1010 260
rect 1010 233 1019 260
rect 967 208 1019 233
rect 1123 1203 1175 1212
rect 1123 1169 1132 1203
rect 1132 1169 1166 1203
rect 1166 1169 1175 1203
rect 1123 1160 1175 1169
rect 1123 1131 1175 1148
rect 1123 1097 1132 1131
rect 1132 1097 1166 1131
rect 1166 1097 1175 1131
rect 1123 1096 1175 1097
rect 1123 1059 1175 1084
rect 1123 1032 1132 1059
rect 1132 1032 1166 1059
rect 1166 1032 1175 1059
rect 1123 987 1175 1020
rect 1123 968 1132 987
rect 1132 968 1166 987
rect 1166 968 1175 987
rect 1123 953 1132 956
rect 1132 953 1166 956
rect 1166 953 1175 956
rect 1123 915 1175 953
rect 1123 904 1132 915
rect 1132 904 1166 915
rect 1166 904 1175 915
rect 1123 881 1132 892
rect 1132 881 1166 892
rect 1166 881 1175 892
rect 1123 843 1175 881
rect 1123 840 1132 843
rect 1132 840 1166 843
rect 1166 840 1175 843
rect 1123 809 1132 828
rect 1132 809 1166 828
rect 1166 809 1175 828
rect 1123 776 1175 809
rect 1123 737 1132 764
rect 1132 737 1166 764
rect 1166 737 1175 764
rect 1123 712 1175 737
rect 1123 699 1175 700
rect 1123 665 1132 699
rect 1132 665 1166 699
rect 1166 665 1175 699
rect 1123 648 1175 665
rect 1123 627 1175 636
rect 1123 593 1132 627
rect 1132 593 1166 627
rect 1166 593 1175 627
rect 1123 584 1175 593
rect 1279 1563 1331 1588
rect 1279 1536 1288 1563
rect 1288 1536 1322 1563
rect 1322 1536 1331 1563
rect 1279 1491 1331 1524
rect 1279 1472 1288 1491
rect 1288 1472 1322 1491
rect 1322 1472 1331 1491
rect 1279 1457 1288 1460
rect 1288 1457 1322 1460
rect 1322 1457 1331 1460
rect 1279 1419 1331 1457
rect 1279 1408 1288 1419
rect 1288 1408 1322 1419
rect 1322 1408 1331 1419
rect 1279 1385 1288 1396
rect 1288 1385 1322 1396
rect 1322 1385 1331 1396
rect 1279 1347 1331 1385
rect 1279 1344 1288 1347
rect 1288 1344 1322 1347
rect 1322 1344 1331 1347
rect 1279 1313 1288 1332
rect 1288 1313 1322 1332
rect 1322 1313 1331 1332
rect 1279 1280 1331 1313
rect 1279 483 1331 516
rect 1279 464 1288 483
rect 1288 464 1322 483
rect 1322 464 1331 483
rect 1279 449 1288 452
rect 1288 449 1322 452
rect 1322 449 1331 452
rect 1279 411 1331 449
rect 1279 400 1288 411
rect 1288 400 1322 411
rect 1322 400 1331 411
rect 1279 377 1288 388
rect 1288 377 1322 388
rect 1322 377 1331 388
rect 1279 339 1331 377
rect 1279 336 1288 339
rect 1288 336 1322 339
rect 1322 336 1331 339
rect 1279 305 1288 324
rect 1288 305 1322 324
rect 1322 305 1331 324
rect 1279 272 1331 305
rect 1279 233 1288 260
rect 1288 233 1322 260
rect 1322 233 1331 260
rect 1279 208 1331 233
rect 1435 1203 1487 1212
rect 1435 1169 1444 1203
rect 1444 1169 1478 1203
rect 1478 1169 1487 1203
rect 1435 1160 1487 1169
rect 1435 1131 1487 1148
rect 1435 1097 1444 1131
rect 1444 1097 1478 1131
rect 1478 1097 1487 1131
rect 1435 1096 1487 1097
rect 1435 1059 1487 1084
rect 1435 1032 1444 1059
rect 1444 1032 1478 1059
rect 1478 1032 1487 1059
rect 1435 987 1487 1020
rect 1435 968 1444 987
rect 1444 968 1478 987
rect 1478 968 1487 987
rect 1435 953 1444 956
rect 1444 953 1478 956
rect 1478 953 1487 956
rect 1435 915 1487 953
rect 1435 904 1444 915
rect 1444 904 1478 915
rect 1478 904 1487 915
rect 1435 881 1444 892
rect 1444 881 1478 892
rect 1478 881 1487 892
rect 1435 843 1487 881
rect 1435 840 1444 843
rect 1444 840 1478 843
rect 1478 840 1487 843
rect 1435 809 1444 828
rect 1444 809 1478 828
rect 1478 809 1487 828
rect 1435 776 1487 809
rect 1435 737 1444 764
rect 1444 737 1478 764
rect 1478 737 1487 764
rect 1435 712 1487 737
rect 1435 699 1487 700
rect 1435 665 1444 699
rect 1444 665 1478 699
rect 1478 665 1487 699
rect 1435 648 1487 665
rect 1435 627 1487 636
rect 1435 593 1444 627
rect 1444 593 1478 627
rect 1478 593 1487 627
rect 1435 584 1487 593
rect 1591 1563 1643 1588
rect 1591 1536 1600 1563
rect 1600 1536 1634 1563
rect 1634 1536 1643 1563
rect 1591 1491 1643 1524
rect 1591 1472 1600 1491
rect 1600 1472 1634 1491
rect 1634 1472 1643 1491
rect 1591 1457 1600 1460
rect 1600 1457 1634 1460
rect 1634 1457 1643 1460
rect 1591 1419 1643 1457
rect 1591 1408 1600 1419
rect 1600 1408 1634 1419
rect 1634 1408 1643 1419
rect 1591 1385 1600 1396
rect 1600 1385 1634 1396
rect 1634 1385 1643 1396
rect 1591 1347 1643 1385
rect 1591 1344 1600 1347
rect 1600 1344 1634 1347
rect 1634 1344 1643 1347
rect 1591 1313 1600 1332
rect 1600 1313 1634 1332
rect 1634 1313 1643 1332
rect 1591 1280 1643 1313
rect 1591 483 1643 516
rect 1591 464 1600 483
rect 1600 464 1634 483
rect 1634 464 1643 483
rect 1591 449 1600 452
rect 1600 449 1634 452
rect 1634 449 1643 452
rect 1591 411 1643 449
rect 1591 400 1600 411
rect 1600 400 1634 411
rect 1634 400 1643 411
rect 1591 377 1600 388
rect 1600 377 1634 388
rect 1634 377 1643 388
rect 1591 339 1643 377
rect 1591 336 1600 339
rect 1600 336 1634 339
rect 1634 336 1643 339
rect 1591 305 1600 324
rect 1600 305 1634 324
rect 1634 305 1643 324
rect 1591 272 1643 305
rect 1591 233 1600 260
rect 1600 233 1634 260
rect 1634 233 1643 260
rect 1591 208 1643 233
rect 1747 1203 1799 1212
rect 1747 1169 1756 1203
rect 1756 1169 1790 1203
rect 1790 1169 1799 1203
rect 1747 1160 1799 1169
rect 1747 1131 1799 1148
rect 1747 1097 1756 1131
rect 1756 1097 1790 1131
rect 1790 1097 1799 1131
rect 1747 1096 1799 1097
rect 1747 1059 1799 1084
rect 1747 1032 1756 1059
rect 1756 1032 1790 1059
rect 1790 1032 1799 1059
rect 1747 987 1799 1020
rect 1747 968 1756 987
rect 1756 968 1790 987
rect 1790 968 1799 987
rect 1747 953 1756 956
rect 1756 953 1790 956
rect 1790 953 1799 956
rect 1747 915 1799 953
rect 1747 904 1756 915
rect 1756 904 1790 915
rect 1790 904 1799 915
rect 1747 881 1756 892
rect 1756 881 1790 892
rect 1790 881 1799 892
rect 1747 843 1799 881
rect 1747 840 1756 843
rect 1756 840 1790 843
rect 1790 840 1799 843
rect 1747 809 1756 828
rect 1756 809 1790 828
rect 1790 809 1799 828
rect 1747 776 1799 809
rect 1747 737 1756 764
rect 1756 737 1790 764
rect 1790 737 1799 764
rect 1747 712 1799 737
rect 1747 699 1799 700
rect 1747 665 1756 699
rect 1756 665 1790 699
rect 1790 665 1799 699
rect 1747 648 1799 665
rect 1747 627 1799 636
rect 1747 593 1756 627
rect 1756 593 1790 627
rect 1790 593 1799 627
rect 1747 584 1799 593
rect 1903 1563 1955 1588
rect 1903 1536 1912 1563
rect 1912 1536 1946 1563
rect 1946 1536 1955 1563
rect 1903 1491 1955 1524
rect 1903 1472 1912 1491
rect 1912 1472 1946 1491
rect 1946 1472 1955 1491
rect 1903 1457 1912 1460
rect 1912 1457 1946 1460
rect 1946 1457 1955 1460
rect 1903 1419 1955 1457
rect 1903 1408 1912 1419
rect 1912 1408 1946 1419
rect 1946 1408 1955 1419
rect 1903 1385 1912 1396
rect 1912 1385 1946 1396
rect 1946 1385 1955 1396
rect 1903 1347 1955 1385
rect 1903 1344 1912 1347
rect 1912 1344 1946 1347
rect 1946 1344 1955 1347
rect 1903 1313 1912 1332
rect 1912 1313 1946 1332
rect 1946 1313 1955 1332
rect 1903 1280 1955 1313
rect 1903 483 1955 516
rect 1903 464 1912 483
rect 1912 464 1946 483
rect 1946 464 1955 483
rect 1903 449 1912 452
rect 1912 449 1946 452
rect 1946 449 1955 452
rect 1903 411 1955 449
rect 1903 400 1912 411
rect 1912 400 1946 411
rect 1946 400 1955 411
rect 1903 377 1912 388
rect 1912 377 1946 388
rect 1946 377 1955 388
rect 1903 339 1955 377
rect 1903 336 1912 339
rect 1912 336 1946 339
rect 1946 336 1955 339
rect 1903 305 1912 324
rect 1912 305 1946 324
rect 1946 305 1955 324
rect 1903 272 1955 305
rect 1903 233 1912 260
rect 1912 233 1946 260
rect 1946 233 1955 260
rect 1903 208 1955 233
<< metal2 >>
rect 14 1588 2284 1594
rect 14 1536 343 1588
rect 395 1536 655 1588
rect 707 1536 967 1588
rect 1019 1536 1279 1588
rect 1331 1536 1591 1588
rect 1643 1536 1903 1588
rect 1955 1536 2284 1588
rect 14 1524 2284 1536
rect 14 1472 343 1524
rect 395 1472 655 1524
rect 707 1472 967 1524
rect 1019 1472 1279 1524
rect 1331 1472 1591 1524
rect 1643 1472 1903 1524
rect 1955 1472 2284 1524
rect 14 1460 2284 1472
rect 14 1408 343 1460
rect 395 1408 655 1460
rect 707 1408 967 1460
rect 1019 1408 1279 1460
rect 1331 1408 1591 1460
rect 1643 1408 1903 1460
rect 1955 1408 2284 1460
rect 14 1396 2284 1408
rect 14 1344 343 1396
rect 395 1344 655 1396
rect 707 1344 967 1396
rect 1019 1344 1279 1396
rect 1331 1344 1591 1396
rect 1643 1344 1903 1396
rect 1955 1344 2284 1396
rect 14 1332 2284 1344
rect 14 1280 343 1332
rect 395 1280 655 1332
rect 707 1280 967 1332
rect 1019 1280 1279 1332
rect 1331 1280 1591 1332
rect 1643 1280 1903 1332
rect 1955 1280 2284 1332
rect 14 1274 2284 1280
rect 14 1212 2284 1218
rect 14 1160 499 1212
rect 551 1160 811 1212
rect 863 1160 1123 1212
rect 1175 1160 1435 1212
rect 1487 1160 1747 1212
rect 1799 1160 2284 1212
rect 14 1148 2284 1160
rect 14 1096 499 1148
rect 551 1096 811 1148
rect 863 1096 1123 1148
rect 1175 1096 1435 1148
rect 1487 1096 1747 1148
rect 1799 1096 2284 1148
rect 14 1084 2284 1096
rect 14 1032 499 1084
rect 551 1032 811 1084
rect 863 1032 1123 1084
rect 1175 1032 1435 1084
rect 1487 1032 1747 1084
rect 1799 1032 2284 1084
rect 14 1020 2284 1032
rect 14 968 499 1020
rect 551 968 811 1020
rect 863 968 1123 1020
rect 1175 968 1435 1020
rect 1487 968 1747 1020
rect 1799 968 2284 1020
rect 14 956 2284 968
rect 14 904 499 956
rect 551 904 811 956
rect 863 904 1123 956
rect 1175 904 1435 956
rect 1487 904 1747 956
rect 1799 904 2284 956
rect 14 892 2284 904
rect 14 840 499 892
rect 551 840 811 892
rect 863 840 1123 892
rect 1175 840 1435 892
rect 1487 840 1747 892
rect 1799 840 2284 892
rect 14 828 2284 840
rect 14 776 499 828
rect 551 776 811 828
rect 863 776 1123 828
rect 1175 776 1435 828
rect 1487 776 1747 828
rect 1799 776 2284 828
rect 14 764 2284 776
rect 14 712 499 764
rect 551 712 811 764
rect 863 712 1123 764
rect 1175 712 1435 764
rect 1487 712 1747 764
rect 1799 712 2284 764
rect 14 700 2284 712
rect 14 648 499 700
rect 551 648 811 700
rect 863 648 1123 700
rect 1175 648 1435 700
rect 1487 648 1747 700
rect 1799 648 2284 700
rect 14 636 2284 648
rect 14 584 499 636
rect 551 584 811 636
rect 863 584 1123 636
rect 1175 584 1435 636
rect 1487 584 1747 636
rect 1799 584 2284 636
rect 14 578 2284 584
rect 14 516 2284 522
rect 14 464 343 516
rect 395 464 655 516
rect 707 464 967 516
rect 1019 464 1279 516
rect 1331 464 1591 516
rect 1643 464 1903 516
rect 1955 464 2284 516
rect 14 452 2284 464
rect 14 400 343 452
rect 395 400 655 452
rect 707 400 967 452
rect 1019 400 1279 452
rect 1331 400 1591 452
rect 1643 400 1903 452
rect 1955 400 2284 452
rect 14 388 2284 400
rect 14 336 343 388
rect 395 336 655 388
rect 707 336 967 388
rect 1019 336 1279 388
rect 1331 336 1591 388
rect 1643 336 1903 388
rect 1955 336 2284 388
rect 14 324 2284 336
rect 14 272 343 324
rect 395 272 655 324
rect 707 272 967 324
rect 1019 272 1279 324
rect 1331 272 1591 324
rect 1643 272 1903 324
rect 1955 272 2284 324
rect 14 260 2284 272
rect 14 208 343 260
rect 395 208 655 260
rect 707 208 967 260
rect 1019 208 1279 260
rect 1331 208 1591 260
rect 1643 208 1903 260
rect 1955 208 2284 260
rect 14 202 2284 208
<< labels >>
flabel metal1 s 1098 85 1195 120 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal2 s 251 1374 287 1535 0 FreeSans 200 90 0 0 SOURCE
port 3 nsew
flabel metal2 s 308 798 349 1034 0 FreeSans 200 90 0 0 DRAIN
port 1 nsew
flabel metal2 s 248 268 290 464 0 FreeSans 200 90 0 0 SOURCE
port 3 nsew
flabel metal1 s 2198 1221 2257 1251 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 41 1231 100 1261 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel comment s 1929 898 1929 898 0 FreeSans 300 0 0 0 S
flabel comment s 1773 898 1773 898 0 FreeSans 300 0 0 0 S
flabel comment s 1773 898 1773 898 0 FreeSans 300 0 0 0 D
flabel comment s 1617 898 1617 898 0 FreeSans 300 0 0 0 S
flabel comment s 1617 898 1617 898 0 FreeSans 300 0 0 0 S
flabel comment s 1461 898 1461 898 0 FreeSans 300 0 0 0 S
flabel comment s 1461 898 1461 898 0 FreeSans 300 0 0 0 D
flabel comment s 1305 898 1305 898 0 FreeSans 300 0 0 0 D
flabel comment s 1305 898 1305 898 0 FreeSans 300 0 0 0 S
flabel comment s 1149 898 1149 898 0 FreeSans 300 0 0 0 S
flabel comment s 1149 898 1149 898 0 FreeSans 300 0 0 0 S
flabel comment s 993 898 993 898 0 FreeSans 300 0 0 0 D
flabel comment s 993 898 993 898 0 FreeSans 300 0 0 0 S
flabel comment s 837 898 837 898 0 FreeSans 300 0 0 0 D
flabel comment s 837 898 837 898 0 FreeSans 300 0 0 0 S
flabel comment s 681 898 681 898 0 FreeSans 300 0 0 0 S
flabel comment s 681 898 681 898 0 FreeSans 300 0 0 0 S
flabel comment s 525 898 525 898 0 FreeSans 300 0 0 0 D
flabel comment s 525 898 525 898 0 FreeSans 300 0 0 0 S
flabel comment s 369 898 369 898 0 FreeSans 300 0 0 0 S
flabel comment s 369 898 369 898 0 FreeSans 300 0 0 0 S
flabel comment s 2002 867 2002 867 0 FreeSans 400 90 0 0 dummy_poly
flabel comment s 283 840 283 840 0 FreeSans 400 90 0 0 dummy_poly
<< properties >>
string GDS_END 8555000
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8486564
string device primitive
<< end >>
