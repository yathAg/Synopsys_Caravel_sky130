magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -36 679 2888 1471
<< pwell >>
rect 2716 25 2818 159
<< psubdiff >>
rect 2742 109 2792 133
rect 2742 75 2750 109
rect 2784 75 2792 109
rect 2742 51 2792 75
<< nsubdiff >>
rect 2742 1339 2792 1363
rect 2742 1305 2750 1339
rect 2784 1305 2792 1339
rect 2742 1281 2792 1305
<< psubdiffcont >>
rect 2750 75 2784 109
<< nsubdiffcont >>
rect 2750 1305 2784 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 2852 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1786 1130 1820 1397
rect 2002 1130 2036 1397
rect 2218 1130 2252 1397
rect 2434 1130 2468 1397
rect 2646 1130 2680 1397
rect 2750 1339 2784 1397
rect 2750 1289 2784 1305
rect 64 724 98 740
rect 64 674 98 690
rect 1354 724 1388 1096
rect 1354 690 1405 724
rect 1354 318 1388 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1786 17 1820 218
rect 2002 17 2036 218
rect 2218 17 2252 218
rect 2434 17 2468 218
rect 2646 17 2680 218
rect 2750 109 2784 125
rect 2750 17 2784 75
rect 0 -17 2852 17
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_16  sky130_sram_1kbyte_1rw1r_32x256_8_contact_16_0
timestamp 1679235063
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_28  sky130_sram_1kbyte_1rw1r_32x256_8_contact_28_0
timestamp 1679235063
transform 1 0 2742 0 1 1281
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_29  sky130_sram_1kbyte_1rw1r_32x256_8_contact_29_0
timestamp 1679235063
transform 1 0 2742 0 1 51
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m24_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_nmos_m24_w2_000_sli_dli_da_p_0
timestamp 1679235063
transform 1 0 54 0 1 51
box -26 -26 2660 456
use sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m24_w2_000_sli_dli_da_p  sky130_sram_1kbyte_1rw1r_32x256_8_pmos_m24_w2_000_sli_dli_da_p_0
timestamp 1679235063
transform 1 0 54 0 1 963
box -59 -56 2693 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
rlabel locali s 1388 707 1388 707 4 Z
rlabel locali s 1426 0 1426 0 4 gnd
rlabel locali s 1426 1414 1426 1414 4 vdd
<< properties >>
string FIXED_BBOX 0 0 2852 1414
string GDS_END 365390
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 361984
<< end >>
