magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 362 163 551 203
rect 1 27 551 163
rect 30 -17 64 27
rect 362 21 551 27
<< scnmos >>
rect 79 53 109 137
rect 259 53 289 137
rect 343 53 373 137
rect 441 47 471 177
<< scpmoshvt >>
rect 79 297 109 381
rect 271 297 301 381
rect 343 297 373 381
rect 441 297 471 497
<< ndiff >>
rect 388 137 441 177
rect 27 106 79 137
rect 27 72 35 106
rect 69 72 79 106
rect 27 53 79 72
rect 109 97 259 137
rect 109 63 119 97
rect 153 63 215 97
rect 249 63 259 97
rect 109 53 259 63
rect 289 111 343 137
rect 289 77 299 111
rect 333 77 343 111
rect 289 53 343 77
rect 373 97 441 137
rect 373 63 393 97
rect 427 63 441 97
rect 373 53 441 63
rect 388 47 441 53
rect 471 135 525 177
rect 471 101 481 135
rect 515 101 525 135
rect 471 47 525 101
<< pdiff >>
rect 388 485 441 497
rect 388 451 396 485
rect 430 451 441 485
rect 388 417 441 451
rect 388 383 396 417
rect 430 383 441 417
rect 388 381 441 383
rect 27 349 79 381
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 341 165 381
rect 109 307 119 341
rect 153 307 165 341
rect 109 297 165 307
rect 219 354 271 381
rect 219 320 227 354
rect 261 320 271 354
rect 219 297 271 320
rect 301 297 343 381
rect 373 297 441 381
rect 471 454 525 497
rect 471 420 481 454
rect 515 420 525 454
rect 471 386 525 420
rect 471 352 481 386
rect 515 352 525 386
rect 471 297 525 352
<< ndiffc >>
rect 35 72 69 106
rect 119 63 153 97
rect 215 63 249 97
rect 299 77 333 111
rect 393 63 427 97
rect 481 101 515 135
<< pdiffc >>
rect 396 451 430 485
rect 396 383 430 417
rect 35 315 69 349
rect 119 307 153 341
rect 227 320 261 354
rect 481 420 515 454
rect 481 352 515 386
<< poly >>
rect 441 497 471 523
rect 169 473 373 483
rect 169 439 185 473
rect 219 453 373 473
rect 219 439 235 453
rect 169 429 235 439
rect 79 381 109 407
rect 271 381 301 407
rect 343 381 373 453
rect 79 265 109 297
rect 271 265 301 297
rect 22 249 109 265
rect 22 215 35 249
rect 69 215 109 249
rect 22 199 109 215
rect 217 249 301 265
rect 217 215 227 249
rect 261 215 301 249
rect 217 199 301 215
rect 79 137 109 199
rect 259 137 289 199
rect 343 137 373 297
rect 441 265 471 297
rect 415 249 471 265
rect 415 215 425 249
rect 459 215 471 249
rect 415 199 471 215
rect 441 177 471 199
rect 79 27 109 53
rect 259 27 289 53
rect 343 27 373 53
rect 441 21 471 47
<< polycont >>
rect 185 439 219 473
rect 35 215 69 249
rect 227 215 261 249
rect 425 215 459 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 18 349 69 527
rect 383 485 439 527
rect 108 473 347 483
rect 108 439 185 473
rect 219 439 347 473
rect 108 417 347 439
rect 383 451 396 485
rect 430 451 439 485
rect 383 417 439 451
rect 383 383 396 417
rect 430 383 439 417
rect 18 315 35 349
rect 18 299 69 315
rect 119 341 153 377
rect 119 265 153 307
rect 198 354 282 383
rect 383 367 439 383
rect 481 454 535 493
rect 515 420 535 454
rect 481 386 535 420
rect 198 320 227 354
rect 261 333 282 354
rect 515 352 535 386
rect 261 320 447 333
rect 198 299 447 320
rect 481 299 535 352
rect 413 265 447 299
rect 18 249 85 265
rect 18 215 35 249
rect 69 215 85 249
rect 119 249 267 265
rect 119 215 227 249
rect 261 215 267 249
rect 119 199 267 215
rect 413 249 459 265
rect 413 215 425 249
rect 413 199 459 215
rect 119 181 169 199
rect 22 147 169 181
rect 413 165 447 199
rect 22 106 84 147
rect 299 131 447 165
rect 501 152 535 299
rect 481 135 535 152
rect 22 72 35 106
rect 69 72 84 106
rect 22 53 84 72
rect 118 97 265 113
rect 118 63 119 97
rect 153 63 215 97
rect 249 63 265 97
rect 118 17 265 63
rect 299 111 333 131
rect 515 101 535 135
rect 299 61 333 77
rect 367 63 393 97
rect 427 63 443 97
rect 481 83 535 101
rect 367 17 443 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 214 425 248 459 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 SLEEP_B
port 2 nsew signal input
flabel locali s 490 357 524 391 0 FreeSans 400 0 0 0 X
port 7 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
rlabel comment s 0 0 0 0 4 lpflow_inputiso1n_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 2347070
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2342164
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 13.800 0.000 
<< end >>
