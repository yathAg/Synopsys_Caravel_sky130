magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect 22 1127 6234 2367
rect 1214 973 6234 1127
rect 4650 972 5163 973
<< pwell >>
rect 19 231 105 905
rect 323 253 5794 905
rect 323 231 694 253
rect 19 145 694 231
rect 2042 145 4115 253
rect 4777 145 5794 253
<< mvnmos >>
rect 405 279 525 879
rect 691 279 811 879
rect 867 279 987 879
rect 1043 279 1163 879
rect 1219 279 1339 879
rect 1395 279 1515 879
rect 1681 279 1801 879
rect 1857 279 1977 879
rect 2033 279 2153 879
rect 2209 279 2329 879
rect 2495 279 2615 879
rect 2671 279 2791 879
rect 2847 279 2967 879
rect 3023 279 3143 879
rect 3199 279 3319 879
rect 3375 279 3495 879
rect 3551 279 3671 879
rect 3727 279 3847 879
rect 3903 279 4023 879
rect 4079 279 4199 879
rect 4255 279 4375 879
rect 4431 279 4551 879
rect 4607 279 4727 879
rect 4783 279 4903 879
rect 4959 279 5079 879
rect 5135 279 5255 879
rect 5311 279 5431 879
rect 5487 279 5607 879
<< mvpmos >>
rect 405 1193 505 2193
rect 691 1193 791 2193
rect 847 1193 947 2193
rect 1003 1193 1103 2193
rect 1159 1193 1259 2193
rect 1425 1193 1525 2193
rect 1581 1193 1681 2193
rect 1737 1193 1837 2193
rect 1893 1193 1993 2193
rect 2049 1193 2149 2193
rect 2205 1193 2305 2193
rect 2361 1193 2461 2193
rect 2517 1193 2617 2193
rect 2673 1193 2773 2193
rect 2829 1193 2929 2193
rect 2985 1193 3085 2193
rect 3141 1193 3241 2193
rect 3297 1193 3417 2193
rect 3473 1193 3593 2193
rect 3649 1193 3769 2193
rect 3825 1193 3945 2193
rect 4001 1193 4121 2193
rect 4177 1193 4297 2193
rect 4353 1193 4473 2193
rect 4529 1193 4649 2193
rect 4815 1193 4915 2193
rect 4971 1193 5071 2193
rect 5127 1193 5227 2193
rect 5283 1193 5383 2193
rect 5439 1193 5539 2193
rect 5595 1193 5695 2193
rect 5751 1193 5851 2193
rect 5907 1193 6007 2193
<< mvndiff >>
rect 349 801 405 879
rect 349 767 360 801
rect 394 767 405 801
rect 349 733 405 767
rect 349 699 360 733
rect 394 699 405 733
rect 349 665 405 699
rect 349 631 360 665
rect 394 631 405 665
rect 349 597 405 631
rect 349 563 360 597
rect 394 563 405 597
rect 349 529 405 563
rect 349 495 360 529
rect 394 495 405 529
rect 349 461 405 495
rect 349 427 360 461
rect 394 427 405 461
rect 349 393 405 427
rect 349 359 360 393
rect 394 359 405 393
rect 349 325 405 359
rect 349 291 360 325
rect 394 291 405 325
rect 349 279 405 291
rect 525 801 578 879
rect 525 767 536 801
rect 570 767 578 801
rect 525 733 578 767
rect 525 699 536 733
rect 570 699 578 733
rect 525 665 578 699
rect 525 631 536 665
rect 570 631 578 665
rect 525 597 578 631
rect 525 563 536 597
rect 570 563 578 597
rect 525 529 578 563
rect 525 495 536 529
rect 570 495 578 529
rect 525 461 578 495
rect 525 427 536 461
rect 570 427 578 461
rect 525 393 578 427
rect 525 359 536 393
rect 570 359 578 393
rect 525 325 578 359
rect 525 291 536 325
rect 570 291 578 325
rect 525 279 578 291
rect 638 801 691 879
rect 638 767 646 801
rect 680 767 691 801
rect 638 733 691 767
rect 638 699 646 733
rect 680 699 691 733
rect 638 665 691 699
rect 638 631 646 665
rect 680 631 691 665
rect 638 597 691 631
rect 638 563 646 597
rect 680 563 691 597
rect 638 529 691 563
rect 638 495 646 529
rect 680 495 691 529
rect 638 461 691 495
rect 638 427 646 461
rect 680 427 691 461
rect 638 393 691 427
rect 638 359 646 393
rect 680 359 691 393
rect 638 325 691 359
rect 638 291 646 325
rect 680 291 691 325
rect 638 279 691 291
rect 811 801 867 879
rect 811 767 822 801
rect 856 767 867 801
rect 811 733 867 767
rect 811 699 822 733
rect 856 699 867 733
rect 811 665 867 699
rect 811 631 822 665
rect 856 631 867 665
rect 811 597 867 631
rect 811 563 822 597
rect 856 563 867 597
rect 811 529 867 563
rect 811 495 822 529
rect 856 495 867 529
rect 811 461 867 495
rect 811 427 822 461
rect 856 427 867 461
rect 811 393 867 427
rect 811 359 822 393
rect 856 359 867 393
rect 811 325 867 359
rect 811 291 822 325
rect 856 291 867 325
rect 811 279 867 291
rect 987 801 1043 879
rect 987 767 998 801
rect 1032 767 1043 801
rect 987 733 1043 767
rect 987 699 998 733
rect 1032 699 1043 733
rect 987 665 1043 699
rect 987 631 998 665
rect 1032 631 1043 665
rect 987 597 1043 631
rect 987 563 998 597
rect 1032 563 1043 597
rect 987 529 1043 563
rect 987 495 998 529
rect 1032 495 1043 529
rect 987 461 1043 495
rect 987 427 998 461
rect 1032 427 1043 461
rect 987 393 1043 427
rect 987 359 998 393
rect 1032 359 1043 393
rect 987 325 1043 359
rect 987 291 998 325
rect 1032 291 1043 325
rect 987 279 1043 291
rect 1163 801 1219 879
rect 1163 767 1174 801
rect 1208 767 1219 801
rect 1163 733 1219 767
rect 1163 699 1174 733
rect 1208 699 1219 733
rect 1163 665 1219 699
rect 1163 631 1174 665
rect 1208 631 1219 665
rect 1163 597 1219 631
rect 1163 563 1174 597
rect 1208 563 1219 597
rect 1163 529 1219 563
rect 1163 495 1174 529
rect 1208 495 1219 529
rect 1163 461 1219 495
rect 1163 427 1174 461
rect 1208 427 1219 461
rect 1163 393 1219 427
rect 1163 359 1174 393
rect 1208 359 1219 393
rect 1163 325 1219 359
rect 1163 291 1174 325
rect 1208 291 1219 325
rect 1163 279 1219 291
rect 1339 801 1395 879
rect 1339 767 1350 801
rect 1384 767 1395 801
rect 1339 733 1395 767
rect 1339 699 1350 733
rect 1384 699 1395 733
rect 1339 665 1395 699
rect 1339 631 1350 665
rect 1384 631 1395 665
rect 1339 597 1395 631
rect 1339 563 1350 597
rect 1384 563 1395 597
rect 1339 529 1395 563
rect 1339 495 1350 529
rect 1384 495 1395 529
rect 1339 461 1395 495
rect 1339 427 1350 461
rect 1384 427 1395 461
rect 1339 393 1395 427
rect 1339 359 1350 393
rect 1384 359 1395 393
rect 1339 325 1395 359
rect 1339 291 1350 325
rect 1384 291 1395 325
rect 1339 279 1395 291
rect 1515 801 1568 879
rect 1515 767 1526 801
rect 1560 767 1568 801
rect 1515 733 1568 767
rect 1515 699 1526 733
rect 1560 699 1568 733
rect 1515 665 1568 699
rect 1515 631 1526 665
rect 1560 631 1568 665
rect 1515 597 1568 631
rect 1515 563 1526 597
rect 1560 563 1568 597
rect 1515 529 1568 563
rect 1515 495 1526 529
rect 1560 495 1568 529
rect 1515 461 1568 495
rect 1515 427 1526 461
rect 1560 427 1568 461
rect 1515 393 1568 427
rect 1515 359 1526 393
rect 1560 359 1568 393
rect 1515 325 1568 359
rect 1515 291 1526 325
rect 1560 291 1568 325
rect 1515 279 1568 291
rect 1628 801 1681 879
rect 1628 767 1636 801
rect 1670 767 1681 801
rect 1628 733 1681 767
rect 1628 699 1636 733
rect 1670 699 1681 733
rect 1628 665 1681 699
rect 1628 631 1636 665
rect 1670 631 1681 665
rect 1628 597 1681 631
rect 1628 563 1636 597
rect 1670 563 1681 597
rect 1628 529 1681 563
rect 1628 495 1636 529
rect 1670 495 1681 529
rect 1628 461 1681 495
rect 1628 427 1636 461
rect 1670 427 1681 461
rect 1628 393 1681 427
rect 1628 359 1636 393
rect 1670 359 1681 393
rect 1628 325 1681 359
rect 1628 291 1636 325
rect 1670 291 1681 325
rect 1628 279 1681 291
rect 1801 801 1857 879
rect 1801 767 1812 801
rect 1846 767 1857 801
rect 1801 733 1857 767
rect 1801 699 1812 733
rect 1846 699 1857 733
rect 1801 665 1857 699
rect 1801 631 1812 665
rect 1846 631 1857 665
rect 1801 597 1857 631
rect 1801 563 1812 597
rect 1846 563 1857 597
rect 1801 529 1857 563
rect 1801 495 1812 529
rect 1846 495 1857 529
rect 1801 461 1857 495
rect 1801 427 1812 461
rect 1846 427 1857 461
rect 1801 393 1857 427
rect 1801 359 1812 393
rect 1846 359 1857 393
rect 1801 325 1857 359
rect 1801 291 1812 325
rect 1846 291 1857 325
rect 1801 279 1857 291
rect 1977 801 2033 879
rect 1977 767 1988 801
rect 2022 767 2033 801
rect 1977 733 2033 767
rect 1977 699 1988 733
rect 2022 699 2033 733
rect 1977 665 2033 699
rect 1977 631 1988 665
rect 2022 631 2033 665
rect 1977 597 2033 631
rect 1977 563 1988 597
rect 2022 563 2033 597
rect 1977 529 2033 563
rect 1977 495 1988 529
rect 2022 495 2033 529
rect 1977 461 2033 495
rect 1977 427 1988 461
rect 2022 427 2033 461
rect 1977 393 2033 427
rect 1977 359 1988 393
rect 2022 359 2033 393
rect 1977 325 2033 359
rect 1977 291 1988 325
rect 2022 291 2033 325
rect 1977 279 2033 291
rect 2153 801 2209 879
rect 2153 767 2164 801
rect 2198 767 2209 801
rect 2153 733 2209 767
rect 2153 699 2164 733
rect 2198 699 2209 733
rect 2153 665 2209 699
rect 2153 631 2164 665
rect 2198 631 2209 665
rect 2153 597 2209 631
rect 2153 563 2164 597
rect 2198 563 2209 597
rect 2153 529 2209 563
rect 2153 495 2164 529
rect 2198 495 2209 529
rect 2153 461 2209 495
rect 2153 427 2164 461
rect 2198 427 2209 461
rect 2153 393 2209 427
rect 2153 359 2164 393
rect 2198 359 2209 393
rect 2153 325 2209 359
rect 2153 291 2164 325
rect 2198 291 2209 325
rect 2153 279 2209 291
rect 2329 801 2382 879
rect 2329 767 2340 801
rect 2374 767 2382 801
rect 2329 733 2382 767
rect 2329 699 2340 733
rect 2374 699 2382 733
rect 2329 665 2382 699
rect 2329 631 2340 665
rect 2374 631 2382 665
rect 2329 597 2382 631
rect 2329 563 2340 597
rect 2374 563 2382 597
rect 2329 529 2382 563
rect 2329 495 2340 529
rect 2374 495 2382 529
rect 2329 461 2382 495
rect 2329 427 2340 461
rect 2374 427 2382 461
rect 2329 393 2382 427
rect 2329 359 2340 393
rect 2374 359 2382 393
rect 2329 325 2382 359
rect 2329 291 2340 325
rect 2374 291 2382 325
rect 2329 279 2382 291
rect 2442 801 2495 879
rect 2442 767 2450 801
rect 2484 767 2495 801
rect 2442 733 2495 767
rect 2442 699 2450 733
rect 2484 699 2495 733
rect 2442 665 2495 699
rect 2442 631 2450 665
rect 2484 631 2495 665
rect 2442 597 2495 631
rect 2442 563 2450 597
rect 2484 563 2495 597
rect 2442 529 2495 563
rect 2442 495 2450 529
rect 2484 495 2495 529
rect 2442 461 2495 495
rect 2442 427 2450 461
rect 2484 427 2495 461
rect 2442 393 2495 427
rect 2442 359 2450 393
rect 2484 359 2495 393
rect 2442 325 2495 359
rect 2442 291 2450 325
rect 2484 291 2495 325
rect 2442 279 2495 291
rect 2615 801 2671 879
rect 2615 767 2626 801
rect 2660 767 2671 801
rect 2615 733 2671 767
rect 2615 699 2626 733
rect 2660 699 2671 733
rect 2615 665 2671 699
rect 2615 631 2626 665
rect 2660 631 2671 665
rect 2615 597 2671 631
rect 2615 563 2626 597
rect 2660 563 2671 597
rect 2615 529 2671 563
rect 2615 495 2626 529
rect 2660 495 2671 529
rect 2615 461 2671 495
rect 2615 427 2626 461
rect 2660 427 2671 461
rect 2615 393 2671 427
rect 2615 359 2626 393
rect 2660 359 2671 393
rect 2615 325 2671 359
rect 2615 291 2626 325
rect 2660 291 2671 325
rect 2615 279 2671 291
rect 2791 801 2847 879
rect 2791 767 2802 801
rect 2836 767 2847 801
rect 2791 733 2847 767
rect 2791 699 2802 733
rect 2836 699 2847 733
rect 2791 665 2847 699
rect 2791 631 2802 665
rect 2836 631 2847 665
rect 2791 597 2847 631
rect 2791 563 2802 597
rect 2836 563 2847 597
rect 2791 529 2847 563
rect 2791 495 2802 529
rect 2836 495 2847 529
rect 2791 461 2847 495
rect 2791 427 2802 461
rect 2836 427 2847 461
rect 2791 393 2847 427
rect 2791 359 2802 393
rect 2836 359 2847 393
rect 2791 325 2847 359
rect 2791 291 2802 325
rect 2836 291 2847 325
rect 2791 279 2847 291
rect 2967 801 3023 879
rect 2967 767 2978 801
rect 3012 767 3023 801
rect 2967 733 3023 767
rect 2967 699 2978 733
rect 3012 699 3023 733
rect 2967 665 3023 699
rect 2967 631 2978 665
rect 3012 631 3023 665
rect 2967 597 3023 631
rect 2967 563 2978 597
rect 3012 563 3023 597
rect 2967 529 3023 563
rect 2967 495 2978 529
rect 3012 495 3023 529
rect 2967 461 3023 495
rect 2967 427 2978 461
rect 3012 427 3023 461
rect 2967 393 3023 427
rect 2967 359 2978 393
rect 3012 359 3023 393
rect 2967 325 3023 359
rect 2967 291 2978 325
rect 3012 291 3023 325
rect 2967 279 3023 291
rect 3143 801 3199 879
rect 3143 767 3154 801
rect 3188 767 3199 801
rect 3143 733 3199 767
rect 3143 699 3154 733
rect 3188 699 3199 733
rect 3143 665 3199 699
rect 3143 631 3154 665
rect 3188 631 3199 665
rect 3143 597 3199 631
rect 3143 563 3154 597
rect 3188 563 3199 597
rect 3143 529 3199 563
rect 3143 495 3154 529
rect 3188 495 3199 529
rect 3143 461 3199 495
rect 3143 427 3154 461
rect 3188 427 3199 461
rect 3143 393 3199 427
rect 3143 359 3154 393
rect 3188 359 3199 393
rect 3143 325 3199 359
rect 3143 291 3154 325
rect 3188 291 3199 325
rect 3143 279 3199 291
rect 3319 801 3375 879
rect 3319 767 3330 801
rect 3364 767 3375 801
rect 3319 733 3375 767
rect 3319 699 3330 733
rect 3364 699 3375 733
rect 3319 665 3375 699
rect 3319 631 3330 665
rect 3364 631 3375 665
rect 3319 597 3375 631
rect 3319 563 3330 597
rect 3364 563 3375 597
rect 3319 529 3375 563
rect 3319 495 3330 529
rect 3364 495 3375 529
rect 3319 461 3375 495
rect 3319 427 3330 461
rect 3364 427 3375 461
rect 3319 393 3375 427
rect 3319 359 3330 393
rect 3364 359 3375 393
rect 3319 325 3375 359
rect 3319 291 3330 325
rect 3364 291 3375 325
rect 3319 279 3375 291
rect 3495 801 3551 879
rect 3495 767 3506 801
rect 3540 767 3551 801
rect 3495 733 3551 767
rect 3495 699 3506 733
rect 3540 699 3551 733
rect 3495 665 3551 699
rect 3495 631 3506 665
rect 3540 631 3551 665
rect 3495 597 3551 631
rect 3495 563 3506 597
rect 3540 563 3551 597
rect 3495 529 3551 563
rect 3495 495 3506 529
rect 3540 495 3551 529
rect 3495 461 3551 495
rect 3495 427 3506 461
rect 3540 427 3551 461
rect 3495 393 3551 427
rect 3495 359 3506 393
rect 3540 359 3551 393
rect 3495 325 3551 359
rect 3495 291 3506 325
rect 3540 291 3551 325
rect 3495 279 3551 291
rect 3671 801 3727 879
rect 3671 767 3682 801
rect 3716 767 3727 801
rect 3671 733 3727 767
rect 3671 699 3682 733
rect 3716 699 3727 733
rect 3671 665 3727 699
rect 3671 631 3682 665
rect 3716 631 3727 665
rect 3671 597 3727 631
rect 3671 563 3682 597
rect 3716 563 3727 597
rect 3671 529 3727 563
rect 3671 495 3682 529
rect 3716 495 3727 529
rect 3671 461 3727 495
rect 3671 427 3682 461
rect 3716 427 3727 461
rect 3671 393 3727 427
rect 3671 359 3682 393
rect 3716 359 3727 393
rect 3671 325 3727 359
rect 3671 291 3682 325
rect 3716 291 3727 325
rect 3671 279 3727 291
rect 3847 801 3903 879
rect 3847 767 3858 801
rect 3892 767 3903 801
rect 3847 733 3903 767
rect 3847 699 3858 733
rect 3892 699 3903 733
rect 3847 665 3903 699
rect 3847 631 3858 665
rect 3892 631 3903 665
rect 3847 597 3903 631
rect 3847 563 3858 597
rect 3892 563 3903 597
rect 3847 529 3903 563
rect 3847 495 3858 529
rect 3892 495 3903 529
rect 3847 461 3903 495
rect 3847 427 3858 461
rect 3892 427 3903 461
rect 3847 393 3903 427
rect 3847 359 3858 393
rect 3892 359 3903 393
rect 3847 325 3903 359
rect 3847 291 3858 325
rect 3892 291 3903 325
rect 3847 279 3903 291
rect 4023 801 4079 879
rect 4023 767 4034 801
rect 4068 767 4079 801
rect 4023 733 4079 767
rect 4023 699 4034 733
rect 4068 699 4079 733
rect 4023 665 4079 699
rect 4023 631 4034 665
rect 4068 631 4079 665
rect 4023 597 4079 631
rect 4023 563 4034 597
rect 4068 563 4079 597
rect 4023 529 4079 563
rect 4023 495 4034 529
rect 4068 495 4079 529
rect 4023 461 4079 495
rect 4023 427 4034 461
rect 4068 427 4079 461
rect 4023 393 4079 427
rect 4023 359 4034 393
rect 4068 359 4079 393
rect 4023 325 4079 359
rect 4023 291 4034 325
rect 4068 291 4079 325
rect 4023 279 4079 291
rect 4199 801 4255 879
rect 4199 767 4210 801
rect 4244 767 4255 801
rect 4199 733 4255 767
rect 4199 699 4210 733
rect 4244 699 4255 733
rect 4199 665 4255 699
rect 4199 631 4210 665
rect 4244 631 4255 665
rect 4199 597 4255 631
rect 4199 563 4210 597
rect 4244 563 4255 597
rect 4199 529 4255 563
rect 4199 495 4210 529
rect 4244 495 4255 529
rect 4199 461 4255 495
rect 4199 427 4210 461
rect 4244 427 4255 461
rect 4199 393 4255 427
rect 4199 359 4210 393
rect 4244 359 4255 393
rect 4199 325 4255 359
rect 4199 291 4210 325
rect 4244 291 4255 325
rect 4199 279 4255 291
rect 4375 801 4431 879
rect 4375 767 4386 801
rect 4420 767 4431 801
rect 4375 733 4431 767
rect 4375 699 4386 733
rect 4420 699 4431 733
rect 4375 665 4431 699
rect 4375 631 4386 665
rect 4420 631 4431 665
rect 4375 597 4431 631
rect 4375 563 4386 597
rect 4420 563 4431 597
rect 4375 529 4431 563
rect 4375 495 4386 529
rect 4420 495 4431 529
rect 4375 461 4431 495
rect 4375 427 4386 461
rect 4420 427 4431 461
rect 4375 393 4431 427
rect 4375 359 4386 393
rect 4420 359 4431 393
rect 4375 325 4431 359
rect 4375 291 4386 325
rect 4420 291 4431 325
rect 4375 279 4431 291
rect 4551 801 4607 879
rect 4551 767 4562 801
rect 4596 767 4607 801
rect 4551 733 4607 767
rect 4551 699 4562 733
rect 4596 699 4607 733
rect 4551 665 4607 699
rect 4551 631 4562 665
rect 4596 631 4607 665
rect 4551 597 4607 631
rect 4551 563 4562 597
rect 4596 563 4607 597
rect 4551 529 4607 563
rect 4551 495 4562 529
rect 4596 495 4607 529
rect 4551 461 4607 495
rect 4551 427 4562 461
rect 4596 427 4607 461
rect 4551 393 4607 427
rect 4551 359 4562 393
rect 4596 359 4607 393
rect 4551 325 4607 359
rect 4551 291 4562 325
rect 4596 291 4607 325
rect 4551 279 4607 291
rect 4727 801 4783 879
rect 4727 767 4738 801
rect 4772 767 4783 801
rect 4727 733 4783 767
rect 4727 699 4738 733
rect 4772 699 4783 733
rect 4727 665 4783 699
rect 4727 631 4738 665
rect 4772 631 4783 665
rect 4727 597 4783 631
rect 4727 563 4738 597
rect 4772 563 4783 597
rect 4727 529 4783 563
rect 4727 495 4738 529
rect 4772 495 4783 529
rect 4727 461 4783 495
rect 4727 427 4738 461
rect 4772 427 4783 461
rect 4727 393 4783 427
rect 4727 359 4738 393
rect 4772 359 4783 393
rect 4727 325 4783 359
rect 4727 291 4738 325
rect 4772 291 4783 325
rect 4727 279 4783 291
rect 4903 801 4959 879
rect 4903 767 4914 801
rect 4948 767 4959 801
rect 4903 733 4959 767
rect 4903 699 4914 733
rect 4948 699 4959 733
rect 4903 665 4959 699
rect 4903 631 4914 665
rect 4948 631 4959 665
rect 4903 597 4959 631
rect 4903 563 4914 597
rect 4948 563 4959 597
rect 4903 529 4959 563
rect 4903 495 4914 529
rect 4948 495 4959 529
rect 4903 461 4959 495
rect 4903 427 4914 461
rect 4948 427 4959 461
rect 4903 393 4959 427
rect 4903 359 4914 393
rect 4948 359 4959 393
rect 4903 325 4959 359
rect 4903 291 4914 325
rect 4948 291 4959 325
rect 4903 279 4959 291
rect 5079 801 5135 879
rect 5079 767 5090 801
rect 5124 767 5135 801
rect 5079 733 5135 767
rect 5079 699 5090 733
rect 5124 699 5135 733
rect 5079 665 5135 699
rect 5079 631 5090 665
rect 5124 631 5135 665
rect 5079 597 5135 631
rect 5079 563 5090 597
rect 5124 563 5135 597
rect 5079 529 5135 563
rect 5079 495 5090 529
rect 5124 495 5135 529
rect 5079 461 5135 495
rect 5079 427 5090 461
rect 5124 427 5135 461
rect 5079 393 5135 427
rect 5079 359 5090 393
rect 5124 359 5135 393
rect 5079 325 5135 359
rect 5079 291 5090 325
rect 5124 291 5135 325
rect 5079 279 5135 291
rect 5255 801 5311 879
rect 5255 767 5266 801
rect 5300 767 5311 801
rect 5255 733 5311 767
rect 5255 699 5266 733
rect 5300 699 5311 733
rect 5255 665 5311 699
rect 5255 631 5266 665
rect 5300 631 5311 665
rect 5255 597 5311 631
rect 5255 563 5266 597
rect 5300 563 5311 597
rect 5255 529 5311 563
rect 5255 495 5266 529
rect 5300 495 5311 529
rect 5255 461 5311 495
rect 5255 427 5266 461
rect 5300 427 5311 461
rect 5255 393 5311 427
rect 5255 359 5266 393
rect 5300 359 5311 393
rect 5255 325 5311 359
rect 5255 291 5266 325
rect 5300 291 5311 325
rect 5255 279 5311 291
rect 5431 801 5487 879
rect 5431 767 5442 801
rect 5476 767 5487 801
rect 5431 733 5487 767
rect 5431 699 5442 733
rect 5476 699 5487 733
rect 5431 665 5487 699
rect 5431 631 5442 665
rect 5476 631 5487 665
rect 5431 597 5487 631
rect 5431 563 5442 597
rect 5476 563 5487 597
rect 5431 529 5487 563
rect 5431 495 5442 529
rect 5476 495 5487 529
rect 5431 461 5487 495
rect 5431 427 5442 461
rect 5476 427 5487 461
rect 5431 393 5487 427
rect 5431 359 5442 393
rect 5476 359 5487 393
rect 5431 325 5487 359
rect 5431 291 5442 325
rect 5476 291 5487 325
rect 5431 279 5487 291
rect 5607 801 5660 879
rect 5607 767 5618 801
rect 5652 767 5660 801
rect 5607 733 5660 767
rect 5607 699 5618 733
rect 5652 699 5660 733
rect 5607 665 5660 699
rect 5607 631 5618 665
rect 5652 631 5660 665
rect 5607 597 5660 631
rect 5607 563 5618 597
rect 5652 563 5660 597
rect 5607 529 5660 563
rect 5607 495 5618 529
rect 5652 495 5660 529
rect 5607 461 5660 495
rect 5607 427 5618 461
rect 5652 427 5660 461
rect 5607 393 5660 427
rect 5607 359 5618 393
rect 5652 359 5660 393
rect 5607 325 5660 359
rect 5607 291 5618 325
rect 5652 291 5660 325
rect 5607 279 5660 291
<< mvpdiff >>
rect 352 2181 405 2193
rect 352 2147 360 2181
rect 394 2147 405 2181
rect 352 2113 405 2147
rect 352 2079 360 2113
rect 394 2079 405 2113
rect 352 2045 405 2079
rect 352 2011 360 2045
rect 394 2011 405 2045
rect 352 1977 405 2011
rect 352 1943 360 1977
rect 394 1943 405 1977
rect 352 1909 405 1943
rect 352 1875 360 1909
rect 394 1875 405 1909
rect 352 1841 405 1875
rect 352 1807 360 1841
rect 394 1807 405 1841
rect 352 1773 405 1807
rect 352 1739 360 1773
rect 394 1739 405 1773
rect 352 1705 405 1739
rect 352 1671 360 1705
rect 394 1671 405 1705
rect 352 1637 405 1671
rect 352 1603 360 1637
rect 394 1603 405 1637
rect 352 1569 405 1603
rect 352 1535 360 1569
rect 394 1535 405 1569
rect 352 1501 405 1535
rect 352 1467 360 1501
rect 394 1467 405 1501
rect 352 1433 405 1467
rect 352 1399 360 1433
rect 394 1399 405 1433
rect 352 1365 405 1399
rect 352 1331 360 1365
rect 394 1331 405 1365
rect 352 1297 405 1331
rect 352 1263 360 1297
rect 394 1263 405 1297
rect 352 1193 405 1263
rect 505 2181 558 2193
rect 505 2147 516 2181
rect 550 2147 558 2181
rect 505 2113 558 2147
rect 505 2079 516 2113
rect 550 2079 558 2113
rect 505 2045 558 2079
rect 505 2011 516 2045
rect 550 2011 558 2045
rect 505 1977 558 2011
rect 505 1943 516 1977
rect 550 1943 558 1977
rect 505 1909 558 1943
rect 505 1875 516 1909
rect 550 1875 558 1909
rect 505 1841 558 1875
rect 505 1807 516 1841
rect 550 1807 558 1841
rect 505 1773 558 1807
rect 505 1739 516 1773
rect 550 1739 558 1773
rect 505 1705 558 1739
rect 505 1671 516 1705
rect 550 1671 558 1705
rect 505 1637 558 1671
rect 505 1603 516 1637
rect 550 1603 558 1637
rect 505 1569 558 1603
rect 505 1535 516 1569
rect 550 1535 558 1569
rect 505 1501 558 1535
rect 505 1467 516 1501
rect 550 1467 558 1501
rect 505 1433 558 1467
rect 505 1399 516 1433
rect 550 1399 558 1433
rect 505 1365 558 1399
rect 505 1331 516 1365
rect 550 1331 558 1365
rect 505 1297 558 1331
rect 505 1263 516 1297
rect 550 1263 558 1297
rect 505 1193 558 1263
rect 638 2181 691 2193
rect 638 2147 646 2181
rect 680 2147 691 2181
rect 638 2113 691 2147
rect 638 2079 646 2113
rect 680 2079 691 2113
rect 638 2045 691 2079
rect 638 2011 646 2045
rect 680 2011 691 2045
rect 638 1977 691 2011
rect 638 1943 646 1977
rect 680 1943 691 1977
rect 638 1909 691 1943
rect 638 1875 646 1909
rect 680 1875 691 1909
rect 638 1841 691 1875
rect 638 1807 646 1841
rect 680 1807 691 1841
rect 638 1773 691 1807
rect 638 1739 646 1773
rect 680 1739 691 1773
rect 638 1705 691 1739
rect 638 1671 646 1705
rect 680 1671 691 1705
rect 638 1637 691 1671
rect 638 1603 646 1637
rect 680 1603 691 1637
rect 638 1569 691 1603
rect 638 1535 646 1569
rect 680 1535 691 1569
rect 638 1501 691 1535
rect 638 1467 646 1501
rect 680 1467 691 1501
rect 638 1433 691 1467
rect 638 1399 646 1433
rect 680 1399 691 1433
rect 638 1365 691 1399
rect 638 1331 646 1365
rect 680 1331 691 1365
rect 638 1297 691 1331
rect 638 1263 646 1297
rect 680 1263 691 1297
rect 638 1193 691 1263
rect 791 2181 847 2193
rect 791 2147 802 2181
rect 836 2147 847 2181
rect 791 2113 847 2147
rect 791 2079 802 2113
rect 836 2079 847 2113
rect 791 2045 847 2079
rect 791 2011 802 2045
rect 836 2011 847 2045
rect 791 1977 847 2011
rect 791 1943 802 1977
rect 836 1943 847 1977
rect 791 1909 847 1943
rect 791 1875 802 1909
rect 836 1875 847 1909
rect 791 1841 847 1875
rect 791 1807 802 1841
rect 836 1807 847 1841
rect 791 1773 847 1807
rect 791 1739 802 1773
rect 836 1739 847 1773
rect 791 1705 847 1739
rect 791 1671 802 1705
rect 836 1671 847 1705
rect 791 1637 847 1671
rect 791 1603 802 1637
rect 836 1603 847 1637
rect 791 1569 847 1603
rect 791 1535 802 1569
rect 836 1535 847 1569
rect 791 1501 847 1535
rect 791 1467 802 1501
rect 836 1467 847 1501
rect 791 1433 847 1467
rect 791 1399 802 1433
rect 836 1399 847 1433
rect 791 1365 847 1399
rect 791 1331 802 1365
rect 836 1331 847 1365
rect 791 1297 847 1331
rect 791 1263 802 1297
rect 836 1263 847 1297
rect 791 1193 847 1263
rect 947 2181 1003 2193
rect 947 2147 958 2181
rect 992 2147 1003 2181
rect 947 2113 1003 2147
rect 947 2079 958 2113
rect 992 2079 1003 2113
rect 947 2045 1003 2079
rect 947 2011 958 2045
rect 992 2011 1003 2045
rect 947 1977 1003 2011
rect 947 1943 958 1977
rect 992 1943 1003 1977
rect 947 1909 1003 1943
rect 947 1875 958 1909
rect 992 1875 1003 1909
rect 947 1841 1003 1875
rect 947 1807 958 1841
rect 992 1807 1003 1841
rect 947 1773 1003 1807
rect 947 1739 958 1773
rect 992 1739 1003 1773
rect 947 1705 1003 1739
rect 947 1671 958 1705
rect 992 1671 1003 1705
rect 947 1637 1003 1671
rect 947 1603 958 1637
rect 992 1603 1003 1637
rect 947 1569 1003 1603
rect 947 1535 958 1569
rect 992 1535 1003 1569
rect 947 1501 1003 1535
rect 947 1467 958 1501
rect 992 1467 1003 1501
rect 947 1433 1003 1467
rect 947 1399 958 1433
rect 992 1399 1003 1433
rect 947 1365 1003 1399
rect 947 1331 958 1365
rect 992 1331 1003 1365
rect 947 1297 1003 1331
rect 947 1263 958 1297
rect 992 1263 1003 1297
rect 947 1193 1003 1263
rect 1103 2181 1159 2193
rect 1103 2147 1114 2181
rect 1148 2147 1159 2181
rect 1103 2113 1159 2147
rect 1103 2079 1114 2113
rect 1148 2079 1159 2113
rect 1103 2045 1159 2079
rect 1103 2011 1114 2045
rect 1148 2011 1159 2045
rect 1103 1977 1159 2011
rect 1103 1943 1114 1977
rect 1148 1943 1159 1977
rect 1103 1909 1159 1943
rect 1103 1875 1114 1909
rect 1148 1875 1159 1909
rect 1103 1841 1159 1875
rect 1103 1807 1114 1841
rect 1148 1807 1159 1841
rect 1103 1773 1159 1807
rect 1103 1739 1114 1773
rect 1148 1739 1159 1773
rect 1103 1705 1159 1739
rect 1103 1671 1114 1705
rect 1148 1671 1159 1705
rect 1103 1637 1159 1671
rect 1103 1603 1114 1637
rect 1148 1603 1159 1637
rect 1103 1569 1159 1603
rect 1103 1535 1114 1569
rect 1148 1535 1159 1569
rect 1103 1501 1159 1535
rect 1103 1467 1114 1501
rect 1148 1467 1159 1501
rect 1103 1433 1159 1467
rect 1103 1399 1114 1433
rect 1148 1399 1159 1433
rect 1103 1365 1159 1399
rect 1103 1331 1114 1365
rect 1148 1331 1159 1365
rect 1103 1297 1159 1331
rect 1103 1263 1114 1297
rect 1148 1263 1159 1297
rect 1103 1193 1159 1263
rect 1259 2181 1312 2193
rect 1259 2147 1270 2181
rect 1304 2147 1312 2181
rect 1259 2113 1312 2147
rect 1259 2079 1270 2113
rect 1304 2079 1312 2113
rect 1259 2045 1312 2079
rect 1259 2011 1270 2045
rect 1304 2011 1312 2045
rect 1259 1977 1312 2011
rect 1259 1943 1270 1977
rect 1304 1943 1312 1977
rect 1259 1909 1312 1943
rect 1259 1875 1270 1909
rect 1304 1875 1312 1909
rect 1259 1841 1312 1875
rect 1259 1807 1270 1841
rect 1304 1807 1312 1841
rect 1259 1773 1312 1807
rect 1259 1739 1270 1773
rect 1304 1739 1312 1773
rect 1259 1705 1312 1739
rect 1259 1671 1270 1705
rect 1304 1671 1312 1705
rect 1259 1637 1312 1671
rect 1259 1603 1270 1637
rect 1304 1603 1312 1637
rect 1259 1569 1312 1603
rect 1259 1535 1270 1569
rect 1304 1535 1312 1569
rect 1259 1501 1312 1535
rect 1259 1467 1270 1501
rect 1304 1467 1312 1501
rect 1259 1433 1312 1467
rect 1259 1399 1270 1433
rect 1304 1399 1312 1433
rect 1259 1365 1312 1399
rect 1259 1331 1270 1365
rect 1304 1331 1312 1365
rect 1259 1297 1312 1331
rect 1259 1263 1270 1297
rect 1304 1263 1312 1297
rect 1259 1193 1312 1263
rect 1372 2181 1425 2193
rect 1372 2147 1380 2181
rect 1414 2147 1425 2181
rect 1372 2113 1425 2147
rect 1372 2079 1380 2113
rect 1414 2079 1425 2113
rect 1372 2045 1425 2079
rect 1372 2011 1380 2045
rect 1414 2011 1425 2045
rect 1372 1977 1425 2011
rect 1372 1943 1380 1977
rect 1414 1943 1425 1977
rect 1372 1909 1425 1943
rect 1372 1875 1380 1909
rect 1414 1875 1425 1909
rect 1372 1841 1425 1875
rect 1372 1807 1380 1841
rect 1414 1807 1425 1841
rect 1372 1773 1425 1807
rect 1372 1739 1380 1773
rect 1414 1739 1425 1773
rect 1372 1705 1425 1739
rect 1372 1671 1380 1705
rect 1414 1671 1425 1705
rect 1372 1637 1425 1671
rect 1372 1603 1380 1637
rect 1414 1603 1425 1637
rect 1372 1569 1425 1603
rect 1372 1535 1380 1569
rect 1414 1535 1425 1569
rect 1372 1501 1425 1535
rect 1372 1467 1380 1501
rect 1414 1467 1425 1501
rect 1372 1433 1425 1467
rect 1372 1399 1380 1433
rect 1414 1399 1425 1433
rect 1372 1365 1425 1399
rect 1372 1331 1380 1365
rect 1414 1331 1425 1365
rect 1372 1297 1425 1331
rect 1372 1263 1380 1297
rect 1414 1263 1425 1297
rect 1372 1193 1425 1263
rect 1525 2181 1581 2193
rect 1525 2147 1536 2181
rect 1570 2147 1581 2181
rect 1525 2113 1581 2147
rect 1525 2079 1536 2113
rect 1570 2079 1581 2113
rect 1525 2045 1581 2079
rect 1525 2011 1536 2045
rect 1570 2011 1581 2045
rect 1525 1977 1581 2011
rect 1525 1943 1536 1977
rect 1570 1943 1581 1977
rect 1525 1909 1581 1943
rect 1525 1875 1536 1909
rect 1570 1875 1581 1909
rect 1525 1841 1581 1875
rect 1525 1807 1536 1841
rect 1570 1807 1581 1841
rect 1525 1773 1581 1807
rect 1525 1739 1536 1773
rect 1570 1739 1581 1773
rect 1525 1705 1581 1739
rect 1525 1671 1536 1705
rect 1570 1671 1581 1705
rect 1525 1637 1581 1671
rect 1525 1603 1536 1637
rect 1570 1603 1581 1637
rect 1525 1569 1581 1603
rect 1525 1535 1536 1569
rect 1570 1535 1581 1569
rect 1525 1501 1581 1535
rect 1525 1467 1536 1501
rect 1570 1467 1581 1501
rect 1525 1433 1581 1467
rect 1525 1399 1536 1433
rect 1570 1399 1581 1433
rect 1525 1365 1581 1399
rect 1525 1331 1536 1365
rect 1570 1331 1581 1365
rect 1525 1297 1581 1331
rect 1525 1263 1536 1297
rect 1570 1263 1581 1297
rect 1525 1193 1581 1263
rect 1681 2181 1737 2193
rect 1681 2147 1692 2181
rect 1726 2147 1737 2181
rect 1681 2113 1737 2147
rect 1681 2079 1692 2113
rect 1726 2079 1737 2113
rect 1681 2045 1737 2079
rect 1681 2011 1692 2045
rect 1726 2011 1737 2045
rect 1681 1977 1737 2011
rect 1681 1943 1692 1977
rect 1726 1943 1737 1977
rect 1681 1909 1737 1943
rect 1681 1875 1692 1909
rect 1726 1875 1737 1909
rect 1681 1841 1737 1875
rect 1681 1807 1692 1841
rect 1726 1807 1737 1841
rect 1681 1773 1737 1807
rect 1681 1739 1692 1773
rect 1726 1739 1737 1773
rect 1681 1705 1737 1739
rect 1681 1671 1692 1705
rect 1726 1671 1737 1705
rect 1681 1637 1737 1671
rect 1681 1603 1692 1637
rect 1726 1603 1737 1637
rect 1681 1569 1737 1603
rect 1681 1535 1692 1569
rect 1726 1535 1737 1569
rect 1681 1501 1737 1535
rect 1681 1467 1692 1501
rect 1726 1467 1737 1501
rect 1681 1433 1737 1467
rect 1681 1399 1692 1433
rect 1726 1399 1737 1433
rect 1681 1365 1737 1399
rect 1681 1331 1692 1365
rect 1726 1331 1737 1365
rect 1681 1297 1737 1331
rect 1681 1263 1692 1297
rect 1726 1263 1737 1297
rect 1681 1193 1737 1263
rect 1837 2181 1893 2193
rect 1837 2147 1848 2181
rect 1882 2147 1893 2181
rect 1837 2113 1893 2147
rect 1837 2079 1848 2113
rect 1882 2079 1893 2113
rect 1837 2045 1893 2079
rect 1837 2011 1848 2045
rect 1882 2011 1893 2045
rect 1837 1977 1893 2011
rect 1837 1943 1848 1977
rect 1882 1943 1893 1977
rect 1837 1909 1893 1943
rect 1837 1875 1848 1909
rect 1882 1875 1893 1909
rect 1837 1841 1893 1875
rect 1837 1807 1848 1841
rect 1882 1807 1893 1841
rect 1837 1773 1893 1807
rect 1837 1739 1848 1773
rect 1882 1739 1893 1773
rect 1837 1705 1893 1739
rect 1837 1671 1848 1705
rect 1882 1671 1893 1705
rect 1837 1637 1893 1671
rect 1837 1603 1848 1637
rect 1882 1603 1893 1637
rect 1837 1569 1893 1603
rect 1837 1535 1848 1569
rect 1882 1535 1893 1569
rect 1837 1501 1893 1535
rect 1837 1467 1848 1501
rect 1882 1467 1893 1501
rect 1837 1433 1893 1467
rect 1837 1399 1848 1433
rect 1882 1399 1893 1433
rect 1837 1365 1893 1399
rect 1837 1331 1848 1365
rect 1882 1331 1893 1365
rect 1837 1297 1893 1331
rect 1837 1263 1848 1297
rect 1882 1263 1893 1297
rect 1837 1193 1893 1263
rect 1993 2181 2049 2193
rect 1993 2147 2004 2181
rect 2038 2147 2049 2181
rect 1993 2113 2049 2147
rect 1993 2079 2004 2113
rect 2038 2079 2049 2113
rect 1993 2045 2049 2079
rect 1993 2011 2004 2045
rect 2038 2011 2049 2045
rect 1993 1977 2049 2011
rect 1993 1943 2004 1977
rect 2038 1943 2049 1977
rect 1993 1909 2049 1943
rect 1993 1875 2004 1909
rect 2038 1875 2049 1909
rect 1993 1841 2049 1875
rect 1993 1807 2004 1841
rect 2038 1807 2049 1841
rect 1993 1773 2049 1807
rect 1993 1739 2004 1773
rect 2038 1739 2049 1773
rect 1993 1705 2049 1739
rect 1993 1671 2004 1705
rect 2038 1671 2049 1705
rect 1993 1637 2049 1671
rect 1993 1603 2004 1637
rect 2038 1603 2049 1637
rect 1993 1569 2049 1603
rect 1993 1535 2004 1569
rect 2038 1535 2049 1569
rect 1993 1501 2049 1535
rect 1993 1467 2004 1501
rect 2038 1467 2049 1501
rect 1993 1433 2049 1467
rect 1993 1399 2004 1433
rect 2038 1399 2049 1433
rect 1993 1365 2049 1399
rect 1993 1331 2004 1365
rect 2038 1331 2049 1365
rect 1993 1297 2049 1331
rect 1993 1263 2004 1297
rect 2038 1263 2049 1297
rect 1993 1193 2049 1263
rect 2149 2181 2205 2193
rect 2149 2147 2160 2181
rect 2194 2147 2205 2181
rect 2149 2113 2205 2147
rect 2149 2079 2160 2113
rect 2194 2079 2205 2113
rect 2149 2045 2205 2079
rect 2149 2011 2160 2045
rect 2194 2011 2205 2045
rect 2149 1977 2205 2011
rect 2149 1943 2160 1977
rect 2194 1943 2205 1977
rect 2149 1909 2205 1943
rect 2149 1875 2160 1909
rect 2194 1875 2205 1909
rect 2149 1841 2205 1875
rect 2149 1807 2160 1841
rect 2194 1807 2205 1841
rect 2149 1773 2205 1807
rect 2149 1739 2160 1773
rect 2194 1739 2205 1773
rect 2149 1705 2205 1739
rect 2149 1671 2160 1705
rect 2194 1671 2205 1705
rect 2149 1637 2205 1671
rect 2149 1603 2160 1637
rect 2194 1603 2205 1637
rect 2149 1569 2205 1603
rect 2149 1535 2160 1569
rect 2194 1535 2205 1569
rect 2149 1501 2205 1535
rect 2149 1467 2160 1501
rect 2194 1467 2205 1501
rect 2149 1433 2205 1467
rect 2149 1399 2160 1433
rect 2194 1399 2205 1433
rect 2149 1365 2205 1399
rect 2149 1331 2160 1365
rect 2194 1331 2205 1365
rect 2149 1297 2205 1331
rect 2149 1263 2160 1297
rect 2194 1263 2205 1297
rect 2149 1193 2205 1263
rect 2305 2181 2361 2193
rect 2305 2147 2316 2181
rect 2350 2147 2361 2181
rect 2305 2113 2361 2147
rect 2305 2079 2316 2113
rect 2350 2079 2361 2113
rect 2305 2045 2361 2079
rect 2305 2011 2316 2045
rect 2350 2011 2361 2045
rect 2305 1977 2361 2011
rect 2305 1943 2316 1977
rect 2350 1943 2361 1977
rect 2305 1909 2361 1943
rect 2305 1875 2316 1909
rect 2350 1875 2361 1909
rect 2305 1841 2361 1875
rect 2305 1807 2316 1841
rect 2350 1807 2361 1841
rect 2305 1773 2361 1807
rect 2305 1739 2316 1773
rect 2350 1739 2361 1773
rect 2305 1705 2361 1739
rect 2305 1671 2316 1705
rect 2350 1671 2361 1705
rect 2305 1637 2361 1671
rect 2305 1603 2316 1637
rect 2350 1603 2361 1637
rect 2305 1569 2361 1603
rect 2305 1535 2316 1569
rect 2350 1535 2361 1569
rect 2305 1501 2361 1535
rect 2305 1467 2316 1501
rect 2350 1467 2361 1501
rect 2305 1433 2361 1467
rect 2305 1399 2316 1433
rect 2350 1399 2361 1433
rect 2305 1365 2361 1399
rect 2305 1331 2316 1365
rect 2350 1331 2361 1365
rect 2305 1297 2361 1331
rect 2305 1263 2316 1297
rect 2350 1263 2361 1297
rect 2305 1193 2361 1263
rect 2461 2181 2517 2193
rect 2461 2147 2472 2181
rect 2506 2147 2517 2181
rect 2461 2113 2517 2147
rect 2461 2079 2472 2113
rect 2506 2079 2517 2113
rect 2461 2045 2517 2079
rect 2461 2011 2472 2045
rect 2506 2011 2517 2045
rect 2461 1977 2517 2011
rect 2461 1943 2472 1977
rect 2506 1943 2517 1977
rect 2461 1909 2517 1943
rect 2461 1875 2472 1909
rect 2506 1875 2517 1909
rect 2461 1841 2517 1875
rect 2461 1807 2472 1841
rect 2506 1807 2517 1841
rect 2461 1773 2517 1807
rect 2461 1739 2472 1773
rect 2506 1739 2517 1773
rect 2461 1705 2517 1739
rect 2461 1671 2472 1705
rect 2506 1671 2517 1705
rect 2461 1637 2517 1671
rect 2461 1603 2472 1637
rect 2506 1603 2517 1637
rect 2461 1569 2517 1603
rect 2461 1535 2472 1569
rect 2506 1535 2517 1569
rect 2461 1501 2517 1535
rect 2461 1467 2472 1501
rect 2506 1467 2517 1501
rect 2461 1433 2517 1467
rect 2461 1399 2472 1433
rect 2506 1399 2517 1433
rect 2461 1365 2517 1399
rect 2461 1331 2472 1365
rect 2506 1331 2517 1365
rect 2461 1297 2517 1331
rect 2461 1263 2472 1297
rect 2506 1263 2517 1297
rect 2461 1193 2517 1263
rect 2617 2181 2673 2193
rect 2617 2147 2628 2181
rect 2662 2147 2673 2181
rect 2617 2113 2673 2147
rect 2617 2079 2628 2113
rect 2662 2079 2673 2113
rect 2617 2045 2673 2079
rect 2617 2011 2628 2045
rect 2662 2011 2673 2045
rect 2617 1977 2673 2011
rect 2617 1943 2628 1977
rect 2662 1943 2673 1977
rect 2617 1909 2673 1943
rect 2617 1875 2628 1909
rect 2662 1875 2673 1909
rect 2617 1841 2673 1875
rect 2617 1807 2628 1841
rect 2662 1807 2673 1841
rect 2617 1773 2673 1807
rect 2617 1739 2628 1773
rect 2662 1739 2673 1773
rect 2617 1705 2673 1739
rect 2617 1671 2628 1705
rect 2662 1671 2673 1705
rect 2617 1637 2673 1671
rect 2617 1603 2628 1637
rect 2662 1603 2673 1637
rect 2617 1569 2673 1603
rect 2617 1535 2628 1569
rect 2662 1535 2673 1569
rect 2617 1501 2673 1535
rect 2617 1467 2628 1501
rect 2662 1467 2673 1501
rect 2617 1433 2673 1467
rect 2617 1399 2628 1433
rect 2662 1399 2673 1433
rect 2617 1365 2673 1399
rect 2617 1331 2628 1365
rect 2662 1331 2673 1365
rect 2617 1297 2673 1331
rect 2617 1263 2628 1297
rect 2662 1263 2673 1297
rect 2617 1193 2673 1263
rect 2773 2181 2829 2193
rect 2773 2147 2784 2181
rect 2818 2147 2829 2181
rect 2773 2113 2829 2147
rect 2773 2079 2784 2113
rect 2818 2079 2829 2113
rect 2773 2045 2829 2079
rect 2773 2011 2784 2045
rect 2818 2011 2829 2045
rect 2773 1977 2829 2011
rect 2773 1943 2784 1977
rect 2818 1943 2829 1977
rect 2773 1909 2829 1943
rect 2773 1875 2784 1909
rect 2818 1875 2829 1909
rect 2773 1841 2829 1875
rect 2773 1807 2784 1841
rect 2818 1807 2829 1841
rect 2773 1773 2829 1807
rect 2773 1739 2784 1773
rect 2818 1739 2829 1773
rect 2773 1705 2829 1739
rect 2773 1671 2784 1705
rect 2818 1671 2829 1705
rect 2773 1637 2829 1671
rect 2773 1603 2784 1637
rect 2818 1603 2829 1637
rect 2773 1569 2829 1603
rect 2773 1535 2784 1569
rect 2818 1535 2829 1569
rect 2773 1501 2829 1535
rect 2773 1467 2784 1501
rect 2818 1467 2829 1501
rect 2773 1433 2829 1467
rect 2773 1399 2784 1433
rect 2818 1399 2829 1433
rect 2773 1365 2829 1399
rect 2773 1331 2784 1365
rect 2818 1331 2829 1365
rect 2773 1297 2829 1331
rect 2773 1263 2784 1297
rect 2818 1263 2829 1297
rect 2773 1193 2829 1263
rect 2929 2181 2985 2193
rect 2929 2147 2940 2181
rect 2974 2147 2985 2181
rect 2929 2113 2985 2147
rect 2929 2079 2940 2113
rect 2974 2079 2985 2113
rect 2929 2045 2985 2079
rect 2929 2011 2940 2045
rect 2974 2011 2985 2045
rect 2929 1977 2985 2011
rect 2929 1943 2940 1977
rect 2974 1943 2985 1977
rect 2929 1909 2985 1943
rect 2929 1875 2940 1909
rect 2974 1875 2985 1909
rect 2929 1841 2985 1875
rect 2929 1807 2940 1841
rect 2974 1807 2985 1841
rect 2929 1773 2985 1807
rect 2929 1739 2940 1773
rect 2974 1739 2985 1773
rect 2929 1705 2985 1739
rect 2929 1671 2940 1705
rect 2974 1671 2985 1705
rect 2929 1637 2985 1671
rect 2929 1603 2940 1637
rect 2974 1603 2985 1637
rect 2929 1569 2985 1603
rect 2929 1535 2940 1569
rect 2974 1535 2985 1569
rect 2929 1501 2985 1535
rect 2929 1467 2940 1501
rect 2974 1467 2985 1501
rect 2929 1433 2985 1467
rect 2929 1399 2940 1433
rect 2974 1399 2985 1433
rect 2929 1365 2985 1399
rect 2929 1331 2940 1365
rect 2974 1331 2985 1365
rect 2929 1297 2985 1331
rect 2929 1263 2940 1297
rect 2974 1263 2985 1297
rect 2929 1193 2985 1263
rect 3085 2181 3141 2193
rect 3085 2147 3096 2181
rect 3130 2147 3141 2181
rect 3085 2113 3141 2147
rect 3085 2079 3096 2113
rect 3130 2079 3141 2113
rect 3085 2045 3141 2079
rect 3085 2011 3096 2045
rect 3130 2011 3141 2045
rect 3085 1977 3141 2011
rect 3085 1943 3096 1977
rect 3130 1943 3141 1977
rect 3085 1909 3141 1943
rect 3085 1875 3096 1909
rect 3130 1875 3141 1909
rect 3085 1841 3141 1875
rect 3085 1807 3096 1841
rect 3130 1807 3141 1841
rect 3085 1773 3141 1807
rect 3085 1739 3096 1773
rect 3130 1739 3141 1773
rect 3085 1705 3141 1739
rect 3085 1671 3096 1705
rect 3130 1671 3141 1705
rect 3085 1637 3141 1671
rect 3085 1603 3096 1637
rect 3130 1603 3141 1637
rect 3085 1569 3141 1603
rect 3085 1535 3096 1569
rect 3130 1535 3141 1569
rect 3085 1501 3141 1535
rect 3085 1467 3096 1501
rect 3130 1467 3141 1501
rect 3085 1433 3141 1467
rect 3085 1399 3096 1433
rect 3130 1399 3141 1433
rect 3085 1365 3141 1399
rect 3085 1331 3096 1365
rect 3130 1331 3141 1365
rect 3085 1297 3141 1331
rect 3085 1263 3096 1297
rect 3130 1263 3141 1297
rect 3085 1193 3141 1263
rect 3241 2181 3297 2193
rect 3241 2147 3252 2181
rect 3286 2147 3297 2181
rect 3241 2113 3297 2147
rect 3241 2079 3252 2113
rect 3286 2079 3297 2113
rect 3241 2045 3297 2079
rect 3241 2011 3252 2045
rect 3286 2011 3297 2045
rect 3241 1977 3297 2011
rect 3241 1943 3252 1977
rect 3286 1943 3297 1977
rect 3241 1909 3297 1943
rect 3241 1875 3252 1909
rect 3286 1875 3297 1909
rect 3241 1841 3297 1875
rect 3241 1807 3252 1841
rect 3286 1807 3297 1841
rect 3241 1773 3297 1807
rect 3241 1739 3252 1773
rect 3286 1739 3297 1773
rect 3241 1705 3297 1739
rect 3241 1671 3252 1705
rect 3286 1671 3297 1705
rect 3241 1637 3297 1671
rect 3241 1603 3252 1637
rect 3286 1603 3297 1637
rect 3241 1569 3297 1603
rect 3241 1535 3252 1569
rect 3286 1535 3297 1569
rect 3241 1501 3297 1535
rect 3241 1467 3252 1501
rect 3286 1467 3297 1501
rect 3241 1433 3297 1467
rect 3241 1399 3252 1433
rect 3286 1399 3297 1433
rect 3241 1365 3297 1399
rect 3241 1331 3252 1365
rect 3286 1331 3297 1365
rect 3241 1297 3297 1331
rect 3241 1263 3252 1297
rect 3286 1263 3297 1297
rect 3241 1193 3297 1263
rect 3417 2181 3473 2193
rect 3417 2147 3428 2181
rect 3462 2147 3473 2181
rect 3417 2113 3473 2147
rect 3417 2079 3428 2113
rect 3462 2079 3473 2113
rect 3417 2045 3473 2079
rect 3417 2011 3428 2045
rect 3462 2011 3473 2045
rect 3417 1977 3473 2011
rect 3417 1943 3428 1977
rect 3462 1943 3473 1977
rect 3417 1909 3473 1943
rect 3417 1875 3428 1909
rect 3462 1875 3473 1909
rect 3417 1841 3473 1875
rect 3417 1807 3428 1841
rect 3462 1807 3473 1841
rect 3417 1773 3473 1807
rect 3417 1739 3428 1773
rect 3462 1739 3473 1773
rect 3417 1705 3473 1739
rect 3417 1671 3428 1705
rect 3462 1671 3473 1705
rect 3417 1637 3473 1671
rect 3417 1603 3428 1637
rect 3462 1603 3473 1637
rect 3417 1569 3473 1603
rect 3417 1535 3428 1569
rect 3462 1535 3473 1569
rect 3417 1501 3473 1535
rect 3417 1467 3428 1501
rect 3462 1467 3473 1501
rect 3417 1433 3473 1467
rect 3417 1399 3428 1433
rect 3462 1399 3473 1433
rect 3417 1365 3473 1399
rect 3417 1331 3428 1365
rect 3462 1331 3473 1365
rect 3417 1297 3473 1331
rect 3417 1263 3428 1297
rect 3462 1263 3473 1297
rect 3417 1193 3473 1263
rect 3593 2181 3649 2193
rect 3593 2147 3604 2181
rect 3638 2147 3649 2181
rect 3593 2113 3649 2147
rect 3593 2079 3604 2113
rect 3638 2079 3649 2113
rect 3593 2045 3649 2079
rect 3593 2011 3604 2045
rect 3638 2011 3649 2045
rect 3593 1977 3649 2011
rect 3593 1943 3604 1977
rect 3638 1943 3649 1977
rect 3593 1909 3649 1943
rect 3593 1875 3604 1909
rect 3638 1875 3649 1909
rect 3593 1841 3649 1875
rect 3593 1807 3604 1841
rect 3638 1807 3649 1841
rect 3593 1773 3649 1807
rect 3593 1739 3604 1773
rect 3638 1739 3649 1773
rect 3593 1705 3649 1739
rect 3593 1671 3604 1705
rect 3638 1671 3649 1705
rect 3593 1637 3649 1671
rect 3593 1603 3604 1637
rect 3638 1603 3649 1637
rect 3593 1569 3649 1603
rect 3593 1535 3604 1569
rect 3638 1535 3649 1569
rect 3593 1501 3649 1535
rect 3593 1467 3604 1501
rect 3638 1467 3649 1501
rect 3593 1433 3649 1467
rect 3593 1399 3604 1433
rect 3638 1399 3649 1433
rect 3593 1365 3649 1399
rect 3593 1331 3604 1365
rect 3638 1331 3649 1365
rect 3593 1297 3649 1331
rect 3593 1263 3604 1297
rect 3638 1263 3649 1297
rect 3593 1193 3649 1263
rect 3769 2181 3825 2193
rect 3769 2147 3780 2181
rect 3814 2147 3825 2181
rect 3769 2113 3825 2147
rect 3769 2079 3780 2113
rect 3814 2079 3825 2113
rect 3769 2045 3825 2079
rect 3769 2011 3780 2045
rect 3814 2011 3825 2045
rect 3769 1977 3825 2011
rect 3769 1943 3780 1977
rect 3814 1943 3825 1977
rect 3769 1909 3825 1943
rect 3769 1875 3780 1909
rect 3814 1875 3825 1909
rect 3769 1841 3825 1875
rect 3769 1807 3780 1841
rect 3814 1807 3825 1841
rect 3769 1773 3825 1807
rect 3769 1739 3780 1773
rect 3814 1739 3825 1773
rect 3769 1705 3825 1739
rect 3769 1671 3780 1705
rect 3814 1671 3825 1705
rect 3769 1637 3825 1671
rect 3769 1603 3780 1637
rect 3814 1603 3825 1637
rect 3769 1569 3825 1603
rect 3769 1535 3780 1569
rect 3814 1535 3825 1569
rect 3769 1501 3825 1535
rect 3769 1467 3780 1501
rect 3814 1467 3825 1501
rect 3769 1433 3825 1467
rect 3769 1399 3780 1433
rect 3814 1399 3825 1433
rect 3769 1365 3825 1399
rect 3769 1331 3780 1365
rect 3814 1331 3825 1365
rect 3769 1297 3825 1331
rect 3769 1263 3780 1297
rect 3814 1263 3825 1297
rect 3769 1193 3825 1263
rect 3945 2181 4001 2193
rect 3945 2147 3956 2181
rect 3990 2147 4001 2181
rect 3945 2113 4001 2147
rect 3945 2079 3956 2113
rect 3990 2079 4001 2113
rect 3945 2045 4001 2079
rect 3945 2011 3956 2045
rect 3990 2011 4001 2045
rect 3945 1977 4001 2011
rect 3945 1943 3956 1977
rect 3990 1943 4001 1977
rect 3945 1909 4001 1943
rect 3945 1875 3956 1909
rect 3990 1875 4001 1909
rect 3945 1841 4001 1875
rect 3945 1807 3956 1841
rect 3990 1807 4001 1841
rect 3945 1773 4001 1807
rect 3945 1739 3956 1773
rect 3990 1739 4001 1773
rect 3945 1705 4001 1739
rect 3945 1671 3956 1705
rect 3990 1671 4001 1705
rect 3945 1637 4001 1671
rect 3945 1603 3956 1637
rect 3990 1603 4001 1637
rect 3945 1569 4001 1603
rect 3945 1535 3956 1569
rect 3990 1535 4001 1569
rect 3945 1501 4001 1535
rect 3945 1467 3956 1501
rect 3990 1467 4001 1501
rect 3945 1433 4001 1467
rect 3945 1399 3956 1433
rect 3990 1399 4001 1433
rect 3945 1365 4001 1399
rect 3945 1331 3956 1365
rect 3990 1331 4001 1365
rect 3945 1297 4001 1331
rect 3945 1263 3956 1297
rect 3990 1263 4001 1297
rect 3945 1193 4001 1263
rect 4121 2181 4177 2193
rect 4121 2147 4132 2181
rect 4166 2147 4177 2181
rect 4121 2113 4177 2147
rect 4121 2079 4132 2113
rect 4166 2079 4177 2113
rect 4121 2045 4177 2079
rect 4121 2011 4132 2045
rect 4166 2011 4177 2045
rect 4121 1977 4177 2011
rect 4121 1943 4132 1977
rect 4166 1943 4177 1977
rect 4121 1909 4177 1943
rect 4121 1875 4132 1909
rect 4166 1875 4177 1909
rect 4121 1841 4177 1875
rect 4121 1807 4132 1841
rect 4166 1807 4177 1841
rect 4121 1773 4177 1807
rect 4121 1739 4132 1773
rect 4166 1739 4177 1773
rect 4121 1705 4177 1739
rect 4121 1671 4132 1705
rect 4166 1671 4177 1705
rect 4121 1637 4177 1671
rect 4121 1603 4132 1637
rect 4166 1603 4177 1637
rect 4121 1569 4177 1603
rect 4121 1535 4132 1569
rect 4166 1535 4177 1569
rect 4121 1501 4177 1535
rect 4121 1467 4132 1501
rect 4166 1467 4177 1501
rect 4121 1433 4177 1467
rect 4121 1399 4132 1433
rect 4166 1399 4177 1433
rect 4121 1365 4177 1399
rect 4121 1331 4132 1365
rect 4166 1331 4177 1365
rect 4121 1297 4177 1331
rect 4121 1263 4132 1297
rect 4166 1263 4177 1297
rect 4121 1193 4177 1263
rect 4297 2181 4353 2193
rect 4297 2147 4308 2181
rect 4342 2147 4353 2181
rect 4297 2113 4353 2147
rect 4297 2079 4308 2113
rect 4342 2079 4353 2113
rect 4297 2045 4353 2079
rect 4297 2011 4308 2045
rect 4342 2011 4353 2045
rect 4297 1977 4353 2011
rect 4297 1943 4308 1977
rect 4342 1943 4353 1977
rect 4297 1909 4353 1943
rect 4297 1875 4308 1909
rect 4342 1875 4353 1909
rect 4297 1841 4353 1875
rect 4297 1807 4308 1841
rect 4342 1807 4353 1841
rect 4297 1773 4353 1807
rect 4297 1739 4308 1773
rect 4342 1739 4353 1773
rect 4297 1705 4353 1739
rect 4297 1671 4308 1705
rect 4342 1671 4353 1705
rect 4297 1637 4353 1671
rect 4297 1603 4308 1637
rect 4342 1603 4353 1637
rect 4297 1569 4353 1603
rect 4297 1535 4308 1569
rect 4342 1535 4353 1569
rect 4297 1501 4353 1535
rect 4297 1467 4308 1501
rect 4342 1467 4353 1501
rect 4297 1433 4353 1467
rect 4297 1399 4308 1433
rect 4342 1399 4353 1433
rect 4297 1365 4353 1399
rect 4297 1331 4308 1365
rect 4342 1331 4353 1365
rect 4297 1297 4353 1331
rect 4297 1263 4308 1297
rect 4342 1263 4353 1297
rect 4297 1193 4353 1263
rect 4473 2181 4529 2193
rect 4473 2147 4484 2181
rect 4518 2147 4529 2181
rect 4473 2113 4529 2147
rect 4473 2079 4484 2113
rect 4518 2079 4529 2113
rect 4473 2045 4529 2079
rect 4473 2011 4484 2045
rect 4518 2011 4529 2045
rect 4473 1977 4529 2011
rect 4473 1943 4484 1977
rect 4518 1943 4529 1977
rect 4473 1909 4529 1943
rect 4473 1875 4484 1909
rect 4518 1875 4529 1909
rect 4473 1841 4529 1875
rect 4473 1807 4484 1841
rect 4518 1807 4529 1841
rect 4473 1773 4529 1807
rect 4473 1739 4484 1773
rect 4518 1739 4529 1773
rect 4473 1705 4529 1739
rect 4473 1671 4484 1705
rect 4518 1671 4529 1705
rect 4473 1637 4529 1671
rect 4473 1603 4484 1637
rect 4518 1603 4529 1637
rect 4473 1569 4529 1603
rect 4473 1535 4484 1569
rect 4518 1535 4529 1569
rect 4473 1501 4529 1535
rect 4473 1467 4484 1501
rect 4518 1467 4529 1501
rect 4473 1433 4529 1467
rect 4473 1399 4484 1433
rect 4518 1399 4529 1433
rect 4473 1365 4529 1399
rect 4473 1331 4484 1365
rect 4518 1331 4529 1365
rect 4473 1297 4529 1331
rect 4473 1263 4484 1297
rect 4518 1263 4529 1297
rect 4473 1193 4529 1263
rect 4649 2181 4702 2193
rect 4649 2147 4660 2181
rect 4694 2147 4702 2181
rect 4649 2113 4702 2147
rect 4649 2079 4660 2113
rect 4694 2079 4702 2113
rect 4649 2045 4702 2079
rect 4649 2011 4660 2045
rect 4694 2011 4702 2045
rect 4649 1977 4702 2011
rect 4649 1943 4660 1977
rect 4694 1943 4702 1977
rect 4649 1909 4702 1943
rect 4649 1875 4660 1909
rect 4694 1875 4702 1909
rect 4649 1841 4702 1875
rect 4649 1807 4660 1841
rect 4694 1807 4702 1841
rect 4649 1773 4702 1807
rect 4649 1739 4660 1773
rect 4694 1739 4702 1773
rect 4649 1705 4702 1739
rect 4649 1671 4660 1705
rect 4694 1671 4702 1705
rect 4649 1637 4702 1671
rect 4649 1603 4660 1637
rect 4694 1603 4702 1637
rect 4649 1569 4702 1603
rect 4649 1535 4660 1569
rect 4694 1535 4702 1569
rect 4649 1501 4702 1535
rect 4649 1467 4660 1501
rect 4694 1467 4702 1501
rect 4649 1433 4702 1467
rect 4649 1399 4660 1433
rect 4694 1399 4702 1433
rect 4649 1365 4702 1399
rect 4649 1331 4660 1365
rect 4694 1331 4702 1365
rect 4649 1297 4702 1331
rect 4649 1263 4660 1297
rect 4694 1263 4702 1297
rect 4649 1193 4702 1263
rect 4762 2181 4815 2193
rect 4762 2147 4770 2181
rect 4804 2147 4815 2181
rect 4762 2113 4815 2147
rect 4762 2079 4770 2113
rect 4804 2079 4815 2113
rect 4762 2045 4815 2079
rect 4762 2011 4770 2045
rect 4804 2011 4815 2045
rect 4762 1977 4815 2011
rect 4762 1943 4770 1977
rect 4804 1943 4815 1977
rect 4762 1909 4815 1943
rect 4762 1875 4770 1909
rect 4804 1875 4815 1909
rect 4762 1841 4815 1875
rect 4762 1807 4770 1841
rect 4804 1807 4815 1841
rect 4762 1773 4815 1807
rect 4762 1739 4770 1773
rect 4804 1739 4815 1773
rect 4762 1705 4815 1739
rect 4762 1671 4770 1705
rect 4804 1671 4815 1705
rect 4762 1637 4815 1671
rect 4762 1603 4770 1637
rect 4804 1603 4815 1637
rect 4762 1569 4815 1603
rect 4762 1535 4770 1569
rect 4804 1535 4815 1569
rect 4762 1501 4815 1535
rect 4762 1467 4770 1501
rect 4804 1467 4815 1501
rect 4762 1433 4815 1467
rect 4762 1399 4770 1433
rect 4804 1399 4815 1433
rect 4762 1365 4815 1399
rect 4762 1331 4770 1365
rect 4804 1331 4815 1365
rect 4762 1297 4815 1331
rect 4762 1263 4770 1297
rect 4804 1263 4815 1297
rect 4762 1193 4815 1263
rect 4915 2181 4971 2193
rect 4915 2147 4926 2181
rect 4960 2147 4971 2181
rect 4915 2113 4971 2147
rect 4915 2079 4926 2113
rect 4960 2079 4971 2113
rect 4915 2045 4971 2079
rect 4915 2011 4926 2045
rect 4960 2011 4971 2045
rect 4915 1977 4971 2011
rect 4915 1943 4926 1977
rect 4960 1943 4971 1977
rect 4915 1909 4971 1943
rect 4915 1875 4926 1909
rect 4960 1875 4971 1909
rect 4915 1841 4971 1875
rect 4915 1807 4926 1841
rect 4960 1807 4971 1841
rect 4915 1773 4971 1807
rect 4915 1739 4926 1773
rect 4960 1739 4971 1773
rect 4915 1705 4971 1739
rect 4915 1671 4926 1705
rect 4960 1671 4971 1705
rect 4915 1637 4971 1671
rect 4915 1603 4926 1637
rect 4960 1603 4971 1637
rect 4915 1569 4971 1603
rect 4915 1535 4926 1569
rect 4960 1535 4971 1569
rect 4915 1501 4971 1535
rect 4915 1467 4926 1501
rect 4960 1467 4971 1501
rect 4915 1433 4971 1467
rect 4915 1399 4926 1433
rect 4960 1399 4971 1433
rect 4915 1365 4971 1399
rect 4915 1331 4926 1365
rect 4960 1331 4971 1365
rect 4915 1297 4971 1331
rect 4915 1263 4926 1297
rect 4960 1263 4971 1297
rect 4915 1193 4971 1263
rect 5071 2181 5127 2193
rect 5071 2147 5082 2181
rect 5116 2147 5127 2181
rect 5071 2113 5127 2147
rect 5071 2079 5082 2113
rect 5116 2079 5127 2113
rect 5071 2045 5127 2079
rect 5071 2011 5082 2045
rect 5116 2011 5127 2045
rect 5071 1977 5127 2011
rect 5071 1943 5082 1977
rect 5116 1943 5127 1977
rect 5071 1909 5127 1943
rect 5071 1875 5082 1909
rect 5116 1875 5127 1909
rect 5071 1841 5127 1875
rect 5071 1807 5082 1841
rect 5116 1807 5127 1841
rect 5071 1773 5127 1807
rect 5071 1739 5082 1773
rect 5116 1739 5127 1773
rect 5071 1705 5127 1739
rect 5071 1671 5082 1705
rect 5116 1671 5127 1705
rect 5071 1637 5127 1671
rect 5071 1603 5082 1637
rect 5116 1603 5127 1637
rect 5071 1569 5127 1603
rect 5071 1535 5082 1569
rect 5116 1535 5127 1569
rect 5071 1501 5127 1535
rect 5071 1467 5082 1501
rect 5116 1467 5127 1501
rect 5071 1433 5127 1467
rect 5071 1399 5082 1433
rect 5116 1399 5127 1433
rect 5071 1365 5127 1399
rect 5071 1331 5082 1365
rect 5116 1331 5127 1365
rect 5071 1297 5127 1331
rect 5071 1263 5082 1297
rect 5116 1263 5127 1297
rect 5071 1193 5127 1263
rect 5227 2181 5283 2193
rect 5227 2147 5238 2181
rect 5272 2147 5283 2181
rect 5227 2113 5283 2147
rect 5227 2079 5238 2113
rect 5272 2079 5283 2113
rect 5227 2045 5283 2079
rect 5227 2011 5238 2045
rect 5272 2011 5283 2045
rect 5227 1977 5283 2011
rect 5227 1943 5238 1977
rect 5272 1943 5283 1977
rect 5227 1909 5283 1943
rect 5227 1875 5238 1909
rect 5272 1875 5283 1909
rect 5227 1841 5283 1875
rect 5227 1807 5238 1841
rect 5272 1807 5283 1841
rect 5227 1773 5283 1807
rect 5227 1739 5238 1773
rect 5272 1739 5283 1773
rect 5227 1705 5283 1739
rect 5227 1671 5238 1705
rect 5272 1671 5283 1705
rect 5227 1637 5283 1671
rect 5227 1603 5238 1637
rect 5272 1603 5283 1637
rect 5227 1569 5283 1603
rect 5227 1535 5238 1569
rect 5272 1535 5283 1569
rect 5227 1501 5283 1535
rect 5227 1467 5238 1501
rect 5272 1467 5283 1501
rect 5227 1433 5283 1467
rect 5227 1399 5238 1433
rect 5272 1399 5283 1433
rect 5227 1365 5283 1399
rect 5227 1331 5238 1365
rect 5272 1331 5283 1365
rect 5227 1297 5283 1331
rect 5227 1263 5238 1297
rect 5272 1263 5283 1297
rect 5227 1193 5283 1263
rect 5383 2181 5439 2193
rect 5383 2147 5394 2181
rect 5428 2147 5439 2181
rect 5383 2113 5439 2147
rect 5383 2079 5394 2113
rect 5428 2079 5439 2113
rect 5383 2045 5439 2079
rect 5383 2011 5394 2045
rect 5428 2011 5439 2045
rect 5383 1977 5439 2011
rect 5383 1943 5394 1977
rect 5428 1943 5439 1977
rect 5383 1909 5439 1943
rect 5383 1875 5394 1909
rect 5428 1875 5439 1909
rect 5383 1841 5439 1875
rect 5383 1807 5394 1841
rect 5428 1807 5439 1841
rect 5383 1773 5439 1807
rect 5383 1739 5394 1773
rect 5428 1739 5439 1773
rect 5383 1705 5439 1739
rect 5383 1671 5394 1705
rect 5428 1671 5439 1705
rect 5383 1637 5439 1671
rect 5383 1603 5394 1637
rect 5428 1603 5439 1637
rect 5383 1569 5439 1603
rect 5383 1535 5394 1569
rect 5428 1535 5439 1569
rect 5383 1501 5439 1535
rect 5383 1467 5394 1501
rect 5428 1467 5439 1501
rect 5383 1433 5439 1467
rect 5383 1399 5394 1433
rect 5428 1399 5439 1433
rect 5383 1365 5439 1399
rect 5383 1331 5394 1365
rect 5428 1331 5439 1365
rect 5383 1297 5439 1331
rect 5383 1263 5394 1297
rect 5428 1263 5439 1297
rect 5383 1193 5439 1263
rect 5539 2181 5595 2193
rect 5539 2147 5550 2181
rect 5584 2147 5595 2181
rect 5539 2113 5595 2147
rect 5539 2079 5550 2113
rect 5584 2079 5595 2113
rect 5539 2045 5595 2079
rect 5539 2011 5550 2045
rect 5584 2011 5595 2045
rect 5539 1977 5595 2011
rect 5539 1943 5550 1977
rect 5584 1943 5595 1977
rect 5539 1909 5595 1943
rect 5539 1875 5550 1909
rect 5584 1875 5595 1909
rect 5539 1841 5595 1875
rect 5539 1807 5550 1841
rect 5584 1807 5595 1841
rect 5539 1773 5595 1807
rect 5539 1739 5550 1773
rect 5584 1739 5595 1773
rect 5539 1705 5595 1739
rect 5539 1671 5550 1705
rect 5584 1671 5595 1705
rect 5539 1637 5595 1671
rect 5539 1603 5550 1637
rect 5584 1603 5595 1637
rect 5539 1569 5595 1603
rect 5539 1535 5550 1569
rect 5584 1535 5595 1569
rect 5539 1501 5595 1535
rect 5539 1467 5550 1501
rect 5584 1467 5595 1501
rect 5539 1433 5595 1467
rect 5539 1399 5550 1433
rect 5584 1399 5595 1433
rect 5539 1365 5595 1399
rect 5539 1331 5550 1365
rect 5584 1331 5595 1365
rect 5539 1297 5595 1331
rect 5539 1263 5550 1297
rect 5584 1263 5595 1297
rect 5539 1193 5595 1263
rect 5695 2181 5751 2193
rect 5695 2147 5706 2181
rect 5740 2147 5751 2181
rect 5695 2113 5751 2147
rect 5695 2079 5706 2113
rect 5740 2079 5751 2113
rect 5695 2045 5751 2079
rect 5695 2011 5706 2045
rect 5740 2011 5751 2045
rect 5695 1977 5751 2011
rect 5695 1943 5706 1977
rect 5740 1943 5751 1977
rect 5695 1909 5751 1943
rect 5695 1875 5706 1909
rect 5740 1875 5751 1909
rect 5695 1841 5751 1875
rect 5695 1807 5706 1841
rect 5740 1807 5751 1841
rect 5695 1773 5751 1807
rect 5695 1739 5706 1773
rect 5740 1739 5751 1773
rect 5695 1705 5751 1739
rect 5695 1671 5706 1705
rect 5740 1671 5751 1705
rect 5695 1637 5751 1671
rect 5695 1603 5706 1637
rect 5740 1603 5751 1637
rect 5695 1569 5751 1603
rect 5695 1535 5706 1569
rect 5740 1535 5751 1569
rect 5695 1501 5751 1535
rect 5695 1467 5706 1501
rect 5740 1467 5751 1501
rect 5695 1433 5751 1467
rect 5695 1399 5706 1433
rect 5740 1399 5751 1433
rect 5695 1365 5751 1399
rect 5695 1331 5706 1365
rect 5740 1331 5751 1365
rect 5695 1297 5751 1331
rect 5695 1263 5706 1297
rect 5740 1263 5751 1297
rect 5695 1193 5751 1263
rect 5851 2181 5907 2193
rect 5851 2147 5862 2181
rect 5896 2147 5907 2181
rect 5851 2113 5907 2147
rect 5851 2079 5862 2113
rect 5896 2079 5907 2113
rect 5851 2045 5907 2079
rect 5851 2011 5862 2045
rect 5896 2011 5907 2045
rect 5851 1977 5907 2011
rect 5851 1943 5862 1977
rect 5896 1943 5907 1977
rect 5851 1909 5907 1943
rect 5851 1875 5862 1909
rect 5896 1875 5907 1909
rect 5851 1841 5907 1875
rect 5851 1807 5862 1841
rect 5896 1807 5907 1841
rect 5851 1773 5907 1807
rect 5851 1739 5862 1773
rect 5896 1739 5907 1773
rect 5851 1705 5907 1739
rect 5851 1671 5862 1705
rect 5896 1671 5907 1705
rect 5851 1637 5907 1671
rect 5851 1603 5862 1637
rect 5896 1603 5907 1637
rect 5851 1569 5907 1603
rect 5851 1535 5862 1569
rect 5896 1535 5907 1569
rect 5851 1501 5907 1535
rect 5851 1467 5862 1501
rect 5896 1467 5907 1501
rect 5851 1433 5907 1467
rect 5851 1399 5862 1433
rect 5896 1399 5907 1433
rect 5851 1365 5907 1399
rect 5851 1331 5862 1365
rect 5896 1331 5907 1365
rect 5851 1297 5907 1331
rect 5851 1263 5862 1297
rect 5896 1263 5907 1297
rect 5851 1193 5907 1263
rect 6007 2181 6060 2193
rect 6007 2147 6018 2181
rect 6052 2147 6060 2181
rect 6007 2113 6060 2147
rect 6007 2079 6018 2113
rect 6052 2079 6060 2113
rect 6007 2045 6060 2079
rect 6007 2011 6018 2045
rect 6052 2011 6060 2045
rect 6007 1977 6060 2011
rect 6007 1943 6018 1977
rect 6052 1943 6060 1977
rect 6007 1909 6060 1943
rect 6007 1875 6018 1909
rect 6052 1875 6060 1909
rect 6007 1841 6060 1875
rect 6007 1807 6018 1841
rect 6052 1807 6060 1841
rect 6007 1773 6060 1807
rect 6007 1739 6018 1773
rect 6052 1739 6060 1773
rect 6007 1705 6060 1739
rect 6007 1671 6018 1705
rect 6052 1671 6060 1705
rect 6007 1637 6060 1671
rect 6007 1603 6018 1637
rect 6052 1603 6060 1637
rect 6007 1569 6060 1603
rect 6007 1535 6018 1569
rect 6052 1535 6060 1569
rect 6007 1501 6060 1535
rect 6007 1467 6018 1501
rect 6052 1467 6060 1501
rect 6007 1433 6060 1467
rect 6007 1399 6018 1433
rect 6052 1399 6060 1433
rect 6007 1365 6060 1399
rect 6007 1331 6018 1365
rect 6052 1331 6060 1365
rect 6007 1297 6060 1331
rect 6007 1263 6018 1297
rect 6052 1263 6060 1297
rect 6007 1193 6060 1263
<< mvndiffc >>
rect 360 767 394 801
rect 360 699 394 733
rect 360 631 394 665
rect 360 563 394 597
rect 360 495 394 529
rect 360 427 394 461
rect 360 359 394 393
rect 360 291 394 325
rect 536 767 570 801
rect 536 699 570 733
rect 536 631 570 665
rect 536 563 570 597
rect 536 495 570 529
rect 536 427 570 461
rect 536 359 570 393
rect 536 291 570 325
rect 646 767 680 801
rect 646 699 680 733
rect 646 631 680 665
rect 646 563 680 597
rect 646 495 680 529
rect 646 427 680 461
rect 646 359 680 393
rect 646 291 680 325
rect 822 767 856 801
rect 822 699 856 733
rect 822 631 856 665
rect 822 563 856 597
rect 822 495 856 529
rect 822 427 856 461
rect 822 359 856 393
rect 822 291 856 325
rect 998 767 1032 801
rect 998 699 1032 733
rect 998 631 1032 665
rect 998 563 1032 597
rect 998 495 1032 529
rect 998 427 1032 461
rect 998 359 1032 393
rect 998 291 1032 325
rect 1174 767 1208 801
rect 1174 699 1208 733
rect 1174 631 1208 665
rect 1174 563 1208 597
rect 1174 495 1208 529
rect 1174 427 1208 461
rect 1174 359 1208 393
rect 1174 291 1208 325
rect 1350 767 1384 801
rect 1350 699 1384 733
rect 1350 631 1384 665
rect 1350 563 1384 597
rect 1350 495 1384 529
rect 1350 427 1384 461
rect 1350 359 1384 393
rect 1350 291 1384 325
rect 1526 767 1560 801
rect 1526 699 1560 733
rect 1526 631 1560 665
rect 1526 563 1560 597
rect 1526 495 1560 529
rect 1526 427 1560 461
rect 1526 359 1560 393
rect 1526 291 1560 325
rect 1636 767 1670 801
rect 1636 699 1670 733
rect 1636 631 1670 665
rect 1636 563 1670 597
rect 1636 495 1670 529
rect 1636 427 1670 461
rect 1636 359 1670 393
rect 1636 291 1670 325
rect 1812 767 1846 801
rect 1812 699 1846 733
rect 1812 631 1846 665
rect 1812 563 1846 597
rect 1812 495 1846 529
rect 1812 427 1846 461
rect 1812 359 1846 393
rect 1812 291 1846 325
rect 1988 767 2022 801
rect 1988 699 2022 733
rect 1988 631 2022 665
rect 1988 563 2022 597
rect 1988 495 2022 529
rect 1988 427 2022 461
rect 1988 359 2022 393
rect 1988 291 2022 325
rect 2164 767 2198 801
rect 2164 699 2198 733
rect 2164 631 2198 665
rect 2164 563 2198 597
rect 2164 495 2198 529
rect 2164 427 2198 461
rect 2164 359 2198 393
rect 2164 291 2198 325
rect 2340 767 2374 801
rect 2340 699 2374 733
rect 2340 631 2374 665
rect 2340 563 2374 597
rect 2340 495 2374 529
rect 2340 427 2374 461
rect 2340 359 2374 393
rect 2340 291 2374 325
rect 2450 767 2484 801
rect 2450 699 2484 733
rect 2450 631 2484 665
rect 2450 563 2484 597
rect 2450 495 2484 529
rect 2450 427 2484 461
rect 2450 359 2484 393
rect 2450 291 2484 325
rect 2626 767 2660 801
rect 2626 699 2660 733
rect 2626 631 2660 665
rect 2626 563 2660 597
rect 2626 495 2660 529
rect 2626 427 2660 461
rect 2626 359 2660 393
rect 2626 291 2660 325
rect 2802 767 2836 801
rect 2802 699 2836 733
rect 2802 631 2836 665
rect 2802 563 2836 597
rect 2802 495 2836 529
rect 2802 427 2836 461
rect 2802 359 2836 393
rect 2802 291 2836 325
rect 2978 767 3012 801
rect 2978 699 3012 733
rect 2978 631 3012 665
rect 2978 563 3012 597
rect 2978 495 3012 529
rect 2978 427 3012 461
rect 2978 359 3012 393
rect 2978 291 3012 325
rect 3154 767 3188 801
rect 3154 699 3188 733
rect 3154 631 3188 665
rect 3154 563 3188 597
rect 3154 495 3188 529
rect 3154 427 3188 461
rect 3154 359 3188 393
rect 3154 291 3188 325
rect 3330 767 3364 801
rect 3330 699 3364 733
rect 3330 631 3364 665
rect 3330 563 3364 597
rect 3330 495 3364 529
rect 3330 427 3364 461
rect 3330 359 3364 393
rect 3330 291 3364 325
rect 3506 767 3540 801
rect 3506 699 3540 733
rect 3506 631 3540 665
rect 3506 563 3540 597
rect 3506 495 3540 529
rect 3506 427 3540 461
rect 3506 359 3540 393
rect 3506 291 3540 325
rect 3682 767 3716 801
rect 3682 699 3716 733
rect 3682 631 3716 665
rect 3682 563 3716 597
rect 3682 495 3716 529
rect 3682 427 3716 461
rect 3682 359 3716 393
rect 3682 291 3716 325
rect 3858 767 3892 801
rect 3858 699 3892 733
rect 3858 631 3892 665
rect 3858 563 3892 597
rect 3858 495 3892 529
rect 3858 427 3892 461
rect 3858 359 3892 393
rect 3858 291 3892 325
rect 4034 767 4068 801
rect 4034 699 4068 733
rect 4034 631 4068 665
rect 4034 563 4068 597
rect 4034 495 4068 529
rect 4034 427 4068 461
rect 4034 359 4068 393
rect 4034 291 4068 325
rect 4210 767 4244 801
rect 4210 699 4244 733
rect 4210 631 4244 665
rect 4210 563 4244 597
rect 4210 495 4244 529
rect 4210 427 4244 461
rect 4210 359 4244 393
rect 4210 291 4244 325
rect 4386 767 4420 801
rect 4386 699 4420 733
rect 4386 631 4420 665
rect 4386 563 4420 597
rect 4386 495 4420 529
rect 4386 427 4420 461
rect 4386 359 4420 393
rect 4386 291 4420 325
rect 4562 767 4596 801
rect 4562 699 4596 733
rect 4562 631 4596 665
rect 4562 563 4596 597
rect 4562 495 4596 529
rect 4562 427 4596 461
rect 4562 359 4596 393
rect 4562 291 4596 325
rect 4738 767 4772 801
rect 4738 699 4772 733
rect 4738 631 4772 665
rect 4738 563 4772 597
rect 4738 495 4772 529
rect 4738 427 4772 461
rect 4738 359 4772 393
rect 4738 291 4772 325
rect 4914 767 4948 801
rect 4914 699 4948 733
rect 4914 631 4948 665
rect 4914 563 4948 597
rect 4914 495 4948 529
rect 4914 427 4948 461
rect 4914 359 4948 393
rect 4914 291 4948 325
rect 5090 767 5124 801
rect 5090 699 5124 733
rect 5090 631 5124 665
rect 5090 563 5124 597
rect 5090 495 5124 529
rect 5090 427 5124 461
rect 5090 359 5124 393
rect 5090 291 5124 325
rect 5266 767 5300 801
rect 5266 699 5300 733
rect 5266 631 5300 665
rect 5266 563 5300 597
rect 5266 495 5300 529
rect 5266 427 5300 461
rect 5266 359 5300 393
rect 5266 291 5300 325
rect 5442 767 5476 801
rect 5442 699 5476 733
rect 5442 631 5476 665
rect 5442 563 5476 597
rect 5442 495 5476 529
rect 5442 427 5476 461
rect 5442 359 5476 393
rect 5442 291 5476 325
rect 5618 767 5652 801
rect 5618 699 5652 733
rect 5618 631 5652 665
rect 5618 563 5652 597
rect 5618 495 5652 529
rect 5618 427 5652 461
rect 5618 359 5652 393
rect 5618 291 5652 325
<< mvpdiffc >>
rect 360 2147 394 2181
rect 360 2079 394 2113
rect 360 2011 394 2045
rect 360 1943 394 1977
rect 360 1875 394 1909
rect 360 1807 394 1841
rect 360 1739 394 1773
rect 360 1671 394 1705
rect 360 1603 394 1637
rect 360 1535 394 1569
rect 360 1467 394 1501
rect 360 1399 394 1433
rect 360 1331 394 1365
rect 360 1263 394 1297
rect 516 2147 550 2181
rect 516 2079 550 2113
rect 516 2011 550 2045
rect 516 1943 550 1977
rect 516 1875 550 1909
rect 516 1807 550 1841
rect 516 1739 550 1773
rect 516 1671 550 1705
rect 516 1603 550 1637
rect 516 1535 550 1569
rect 516 1467 550 1501
rect 516 1399 550 1433
rect 516 1331 550 1365
rect 516 1263 550 1297
rect 646 2147 680 2181
rect 646 2079 680 2113
rect 646 2011 680 2045
rect 646 1943 680 1977
rect 646 1875 680 1909
rect 646 1807 680 1841
rect 646 1739 680 1773
rect 646 1671 680 1705
rect 646 1603 680 1637
rect 646 1535 680 1569
rect 646 1467 680 1501
rect 646 1399 680 1433
rect 646 1331 680 1365
rect 646 1263 680 1297
rect 802 2147 836 2181
rect 802 2079 836 2113
rect 802 2011 836 2045
rect 802 1943 836 1977
rect 802 1875 836 1909
rect 802 1807 836 1841
rect 802 1739 836 1773
rect 802 1671 836 1705
rect 802 1603 836 1637
rect 802 1535 836 1569
rect 802 1467 836 1501
rect 802 1399 836 1433
rect 802 1331 836 1365
rect 802 1263 836 1297
rect 958 2147 992 2181
rect 958 2079 992 2113
rect 958 2011 992 2045
rect 958 1943 992 1977
rect 958 1875 992 1909
rect 958 1807 992 1841
rect 958 1739 992 1773
rect 958 1671 992 1705
rect 958 1603 992 1637
rect 958 1535 992 1569
rect 958 1467 992 1501
rect 958 1399 992 1433
rect 958 1331 992 1365
rect 958 1263 992 1297
rect 1114 2147 1148 2181
rect 1114 2079 1148 2113
rect 1114 2011 1148 2045
rect 1114 1943 1148 1977
rect 1114 1875 1148 1909
rect 1114 1807 1148 1841
rect 1114 1739 1148 1773
rect 1114 1671 1148 1705
rect 1114 1603 1148 1637
rect 1114 1535 1148 1569
rect 1114 1467 1148 1501
rect 1114 1399 1148 1433
rect 1114 1331 1148 1365
rect 1114 1263 1148 1297
rect 1270 2147 1304 2181
rect 1270 2079 1304 2113
rect 1270 2011 1304 2045
rect 1270 1943 1304 1977
rect 1270 1875 1304 1909
rect 1270 1807 1304 1841
rect 1270 1739 1304 1773
rect 1270 1671 1304 1705
rect 1270 1603 1304 1637
rect 1270 1535 1304 1569
rect 1270 1467 1304 1501
rect 1270 1399 1304 1433
rect 1270 1331 1304 1365
rect 1270 1263 1304 1297
rect 1380 2147 1414 2181
rect 1380 2079 1414 2113
rect 1380 2011 1414 2045
rect 1380 1943 1414 1977
rect 1380 1875 1414 1909
rect 1380 1807 1414 1841
rect 1380 1739 1414 1773
rect 1380 1671 1414 1705
rect 1380 1603 1414 1637
rect 1380 1535 1414 1569
rect 1380 1467 1414 1501
rect 1380 1399 1414 1433
rect 1380 1331 1414 1365
rect 1380 1263 1414 1297
rect 1536 2147 1570 2181
rect 1536 2079 1570 2113
rect 1536 2011 1570 2045
rect 1536 1943 1570 1977
rect 1536 1875 1570 1909
rect 1536 1807 1570 1841
rect 1536 1739 1570 1773
rect 1536 1671 1570 1705
rect 1536 1603 1570 1637
rect 1536 1535 1570 1569
rect 1536 1467 1570 1501
rect 1536 1399 1570 1433
rect 1536 1331 1570 1365
rect 1536 1263 1570 1297
rect 1692 2147 1726 2181
rect 1692 2079 1726 2113
rect 1692 2011 1726 2045
rect 1692 1943 1726 1977
rect 1692 1875 1726 1909
rect 1692 1807 1726 1841
rect 1692 1739 1726 1773
rect 1692 1671 1726 1705
rect 1692 1603 1726 1637
rect 1692 1535 1726 1569
rect 1692 1467 1726 1501
rect 1692 1399 1726 1433
rect 1692 1331 1726 1365
rect 1692 1263 1726 1297
rect 1848 2147 1882 2181
rect 1848 2079 1882 2113
rect 1848 2011 1882 2045
rect 1848 1943 1882 1977
rect 1848 1875 1882 1909
rect 1848 1807 1882 1841
rect 1848 1739 1882 1773
rect 1848 1671 1882 1705
rect 1848 1603 1882 1637
rect 1848 1535 1882 1569
rect 1848 1467 1882 1501
rect 1848 1399 1882 1433
rect 1848 1331 1882 1365
rect 1848 1263 1882 1297
rect 2004 2147 2038 2181
rect 2004 2079 2038 2113
rect 2004 2011 2038 2045
rect 2004 1943 2038 1977
rect 2004 1875 2038 1909
rect 2004 1807 2038 1841
rect 2004 1739 2038 1773
rect 2004 1671 2038 1705
rect 2004 1603 2038 1637
rect 2004 1535 2038 1569
rect 2004 1467 2038 1501
rect 2004 1399 2038 1433
rect 2004 1331 2038 1365
rect 2004 1263 2038 1297
rect 2160 2147 2194 2181
rect 2160 2079 2194 2113
rect 2160 2011 2194 2045
rect 2160 1943 2194 1977
rect 2160 1875 2194 1909
rect 2160 1807 2194 1841
rect 2160 1739 2194 1773
rect 2160 1671 2194 1705
rect 2160 1603 2194 1637
rect 2160 1535 2194 1569
rect 2160 1467 2194 1501
rect 2160 1399 2194 1433
rect 2160 1331 2194 1365
rect 2160 1263 2194 1297
rect 2316 2147 2350 2181
rect 2316 2079 2350 2113
rect 2316 2011 2350 2045
rect 2316 1943 2350 1977
rect 2316 1875 2350 1909
rect 2316 1807 2350 1841
rect 2316 1739 2350 1773
rect 2316 1671 2350 1705
rect 2316 1603 2350 1637
rect 2316 1535 2350 1569
rect 2316 1467 2350 1501
rect 2316 1399 2350 1433
rect 2316 1331 2350 1365
rect 2316 1263 2350 1297
rect 2472 2147 2506 2181
rect 2472 2079 2506 2113
rect 2472 2011 2506 2045
rect 2472 1943 2506 1977
rect 2472 1875 2506 1909
rect 2472 1807 2506 1841
rect 2472 1739 2506 1773
rect 2472 1671 2506 1705
rect 2472 1603 2506 1637
rect 2472 1535 2506 1569
rect 2472 1467 2506 1501
rect 2472 1399 2506 1433
rect 2472 1331 2506 1365
rect 2472 1263 2506 1297
rect 2628 2147 2662 2181
rect 2628 2079 2662 2113
rect 2628 2011 2662 2045
rect 2628 1943 2662 1977
rect 2628 1875 2662 1909
rect 2628 1807 2662 1841
rect 2628 1739 2662 1773
rect 2628 1671 2662 1705
rect 2628 1603 2662 1637
rect 2628 1535 2662 1569
rect 2628 1467 2662 1501
rect 2628 1399 2662 1433
rect 2628 1331 2662 1365
rect 2628 1263 2662 1297
rect 2784 2147 2818 2181
rect 2784 2079 2818 2113
rect 2784 2011 2818 2045
rect 2784 1943 2818 1977
rect 2784 1875 2818 1909
rect 2784 1807 2818 1841
rect 2784 1739 2818 1773
rect 2784 1671 2818 1705
rect 2784 1603 2818 1637
rect 2784 1535 2818 1569
rect 2784 1467 2818 1501
rect 2784 1399 2818 1433
rect 2784 1331 2818 1365
rect 2784 1263 2818 1297
rect 2940 2147 2974 2181
rect 2940 2079 2974 2113
rect 2940 2011 2974 2045
rect 2940 1943 2974 1977
rect 2940 1875 2974 1909
rect 2940 1807 2974 1841
rect 2940 1739 2974 1773
rect 2940 1671 2974 1705
rect 2940 1603 2974 1637
rect 2940 1535 2974 1569
rect 2940 1467 2974 1501
rect 2940 1399 2974 1433
rect 2940 1331 2974 1365
rect 2940 1263 2974 1297
rect 3096 2147 3130 2181
rect 3096 2079 3130 2113
rect 3096 2011 3130 2045
rect 3096 1943 3130 1977
rect 3096 1875 3130 1909
rect 3096 1807 3130 1841
rect 3096 1739 3130 1773
rect 3096 1671 3130 1705
rect 3096 1603 3130 1637
rect 3096 1535 3130 1569
rect 3096 1467 3130 1501
rect 3096 1399 3130 1433
rect 3096 1331 3130 1365
rect 3096 1263 3130 1297
rect 3252 2147 3286 2181
rect 3252 2079 3286 2113
rect 3252 2011 3286 2045
rect 3252 1943 3286 1977
rect 3252 1875 3286 1909
rect 3252 1807 3286 1841
rect 3252 1739 3286 1773
rect 3252 1671 3286 1705
rect 3252 1603 3286 1637
rect 3252 1535 3286 1569
rect 3252 1467 3286 1501
rect 3252 1399 3286 1433
rect 3252 1331 3286 1365
rect 3252 1263 3286 1297
rect 3428 2147 3462 2181
rect 3428 2079 3462 2113
rect 3428 2011 3462 2045
rect 3428 1943 3462 1977
rect 3428 1875 3462 1909
rect 3428 1807 3462 1841
rect 3428 1739 3462 1773
rect 3428 1671 3462 1705
rect 3428 1603 3462 1637
rect 3428 1535 3462 1569
rect 3428 1467 3462 1501
rect 3428 1399 3462 1433
rect 3428 1331 3462 1365
rect 3428 1263 3462 1297
rect 3604 2147 3638 2181
rect 3604 2079 3638 2113
rect 3604 2011 3638 2045
rect 3604 1943 3638 1977
rect 3604 1875 3638 1909
rect 3604 1807 3638 1841
rect 3604 1739 3638 1773
rect 3604 1671 3638 1705
rect 3604 1603 3638 1637
rect 3604 1535 3638 1569
rect 3604 1467 3638 1501
rect 3604 1399 3638 1433
rect 3604 1331 3638 1365
rect 3604 1263 3638 1297
rect 3780 2147 3814 2181
rect 3780 2079 3814 2113
rect 3780 2011 3814 2045
rect 3780 1943 3814 1977
rect 3780 1875 3814 1909
rect 3780 1807 3814 1841
rect 3780 1739 3814 1773
rect 3780 1671 3814 1705
rect 3780 1603 3814 1637
rect 3780 1535 3814 1569
rect 3780 1467 3814 1501
rect 3780 1399 3814 1433
rect 3780 1331 3814 1365
rect 3780 1263 3814 1297
rect 3956 2147 3990 2181
rect 3956 2079 3990 2113
rect 3956 2011 3990 2045
rect 3956 1943 3990 1977
rect 3956 1875 3990 1909
rect 3956 1807 3990 1841
rect 3956 1739 3990 1773
rect 3956 1671 3990 1705
rect 3956 1603 3990 1637
rect 3956 1535 3990 1569
rect 3956 1467 3990 1501
rect 3956 1399 3990 1433
rect 3956 1331 3990 1365
rect 3956 1263 3990 1297
rect 4132 2147 4166 2181
rect 4132 2079 4166 2113
rect 4132 2011 4166 2045
rect 4132 1943 4166 1977
rect 4132 1875 4166 1909
rect 4132 1807 4166 1841
rect 4132 1739 4166 1773
rect 4132 1671 4166 1705
rect 4132 1603 4166 1637
rect 4132 1535 4166 1569
rect 4132 1467 4166 1501
rect 4132 1399 4166 1433
rect 4132 1331 4166 1365
rect 4132 1263 4166 1297
rect 4308 2147 4342 2181
rect 4308 2079 4342 2113
rect 4308 2011 4342 2045
rect 4308 1943 4342 1977
rect 4308 1875 4342 1909
rect 4308 1807 4342 1841
rect 4308 1739 4342 1773
rect 4308 1671 4342 1705
rect 4308 1603 4342 1637
rect 4308 1535 4342 1569
rect 4308 1467 4342 1501
rect 4308 1399 4342 1433
rect 4308 1331 4342 1365
rect 4308 1263 4342 1297
rect 4484 2147 4518 2181
rect 4484 2079 4518 2113
rect 4484 2011 4518 2045
rect 4484 1943 4518 1977
rect 4484 1875 4518 1909
rect 4484 1807 4518 1841
rect 4484 1739 4518 1773
rect 4484 1671 4518 1705
rect 4484 1603 4518 1637
rect 4484 1535 4518 1569
rect 4484 1467 4518 1501
rect 4484 1399 4518 1433
rect 4484 1331 4518 1365
rect 4484 1263 4518 1297
rect 4660 2147 4694 2181
rect 4660 2079 4694 2113
rect 4660 2011 4694 2045
rect 4660 1943 4694 1977
rect 4660 1875 4694 1909
rect 4660 1807 4694 1841
rect 4660 1739 4694 1773
rect 4660 1671 4694 1705
rect 4660 1603 4694 1637
rect 4660 1535 4694 1569
rect 4660 1467 4694 1501
rect 4660 1399 4694 1433
rect 4660 1331 4694 1365
rect 4660 1263 4694 1297
rect 4770 2147 4804 2181
rect 4770 2079 4804 2113
rect 4770 2011 4804 2045
rect 4770 1943 4804 1977
rect 4770 1875 4804 1909
rect 4770 1807 4804 1841
rect 4770 1739 4804 1773
rect 4770 1671 4804 1705
rect 4770 1603 4804 1637
rect 4770 1535 4804 1569
rect 4770 1467 4804 1501
rect 4770 1399 4804 1433
rect 4770 1331 4804 1365
rect 4770 1263 4804 1297
rect 4926 2147 4960 2181
rect 4926 2079 4960 2113
rect 4926 2011 4960 2045
rect 4926 1943 4960 1977
rect 4926 1875 4960 1909
rect 4926 1807 4960 1841
rect 4926 1739 4960 1773
rect 4926 1671 4960 1705
rect 4926 1603 4960 1637
rect 4926 1535 4960 1569
rect 4926 1467 4960 1501
rect 4926 1399 4960 1433
rect 4926 1331 4960 1365
rect 4926 1263 4960 1297
rect 5082 2147 5116 2181
rect 5082 2079 5116 2113
rect 5082 2011 5116 2045
rect 5082 1943 5116 1977
rect 5082 1875 5116 1909
rect 5082 1807 5116 1841
rect 5082 1739 5116 1773
rect 5082 1671 5116 1705
rect 5082 1603 5116 1637
rect 5082 1535 5116 1569
rect 5082 1467 5116 1501
rect 5082 1399 5116 1433
rect 5082 1331 5116 1365
rect 5082 1263 5116 1297
rect 5238 2147 5272 2181
rect 5238 2079 5272 2113
rect 5238 2011 5272 2045
rect 5238 1943 5272 1977
rect 5238 1875 5272 1909
rect 5238 1807 5272 1841
rect 5238 1739 5272 1773
rect 5238 1671 5272 1705
rect 5238 1603 5272 1637
rect 5238 1535 5272 1569
rect 5238 1467 5272 1501
rect 5238 1399 5272 1433
rect 5238 1331 5272 1365
rect 5238 1263 5272 1297
rect 5394 2147 5428 2181
rect 5394 2079 5428 2113
rect 5394 2011 5428 2045
rect 5394 1943 5428 1977
rect 5394 1875 5428 1909
rect 5394 1807 5428 1841
rect 5394 1739 5428 1773
rect 5394 1671 5428 1705
rect 5394 1603 5428 1637
rect 5394 1535 5428 1569
rect 5394 1467 5428 1501
rect 5394 1399 5428 1433
rect 5394 1331 5428 1365
rect 5394 1263 5428 1297
rect 5550 2147 5584 2181
rect 5550 2079 5584 2113
rect 5550 2011 5584 2045
rect 5550 1943 5584 1977
rect 5550 1875 5584 1909
rect 5550 1807 5584 1841
rect 5550 1739 5584 1773
rect 5550 1671 5584 1705
rect 5550 1603 5584 1637
rect 5550 1535 5584 1569
rect 5550 1467 5584 1501
rect 5550 1399 5584 1433
rect 5550 1331 5584 1365
rect 5550 1263 5584 1297
rect 5706 2147 5740 2181
rect 5706 2079 5740 2113
rect 5706 2011 5740 2045
rect 5706 1943 5740 1977
rect 5706 1875 5740 1909
rect 5706 1807 5740 1841
rect 5706 1739 5740 1773
rect 5706 1671 5740 1705
rect 5706 1603 5740 1637
rect 5706 1535 5740 1569
rect 5706 1467 5740 1501
rect 5706 1399 5740 1433
rect 5706 1331 5740 1365
rect 5706 1263 5740 1297
rect 5862 2147 5896 2181
rect 5862 2079 5896 2113
rect 5862 2011 5896 2045
rect 5862 1943 5896 1977
rect 5862 1875 5896 1909
rect 5862 1807 5896 1841
rect 5862 1739 5896 1773
rect 5862 1671 5896 1705
rect 5862 1603 5896 1637
rect 5862 1535 5896 1569
rect 5862 1467 5896 1501
rect 5862 1399 5896 1433
rect 5862 1331 5896 1365
rect 5862 1263 5896 1297
rect 6018 2147 6052 2181
rect 6018 2079 6052 2113
rect 6018 2011 6052 2045
rect 6018 1943 6052 1977
rect 6018 1875 6052 1909
rect 6018 1807 6052 1841
rect 6018 1739 6052 1773
rect 6018 1671 6052 1705
rect 6018 1603 6052 1637
rect 6018 1535 6052 1569
rect 6018 1467 6052 1501
rect 6018 1399 6052 1433
rect 6018 1331 6052 1365
rect 6018 1263 6052 1297
<< psubdiff >>
rect 45 855 79 879
rect 45 785 79 821
rect 45 715 79 751
rect 45 645 79 681
rect 45 575 79 611
rect 45 506 79 541
rect 45 437 79 472
rect 45 368 79 403
rect 45 299 79 334
rect 5734 855 5768 879
rect 5734 781 5768 821
rect 5734 707 5768 747
rect 5734 633 5768 673
rect 5734 559 5768 599
rect 5734 485 5768 525
rect 5734 411 5768 451
rect 5734 337 5768 377
rect 45 205 79 265
rect 5734 205 5768 303
rect 45 171 69 205
rect 103 171 147 205
rect 181 171 225 205
rect 259 171 302 205
rect 336 171 379 205
rect 413 171 456 205
rect 490 171 533 205
rect 567 171 610 205
rect 644 171 668 205
rect 2068 171 2092 205
rect 2126 171 2162 205
rect 2196 171 2232 205
rect 2266 171 2302 205
rect 2336 171 2372 205
rect 2406 171 2442 205
rect 2476 171 2512 205
rect 2546 171 2582 205
rect 2616 171 2651 205
rect 2685 171 2720 205
rect 2754 171 2789 205
rect 2823 171 2858 205
rect 2892 171 2927 205
rect 2961 171 2996 205
rect 3030 171 3065 205
rect 3099 171 3134 205
rect 3168 171 3203 205
rect 3237 171 3272 205
rect 3306 171 3341 205
rect 3375 171 3410 205
rect 3444 171 3479 205
rect 3513 171 3548 205
rect 3582 171 3617 205
rect 3651 171 3686 205
rect 3720 171 3755 205
rect 3789 171 3824 205
rect 3858 171 3893 205
rect 3927 171 3962 205
rect 3996 171 4031 205
rect 4065 171 4089 205
rect 4803 171 4827 205
rect 4861 171 4901 205
rect 4935 171 4975 205
rect 5009 171 5049 205
rect 5083 171 5123 205
rect 5157 171 5197 205
rect 5231 171 5271 205
rect 5305 171 5345 205
rect 5379 171 5418 205
rect 5452 171 5491 205
rect 5525 171 5564 205
rect 5598 171 5637 205
rect 5671 171 5710 205
rect 5744 171 5768 205
<< mvnsubdiff >>
rect 88 2267 112 2301
rect 146 2267 181 2301
rect 215 2267 250 2301
rect 284 2267 319 2301
rect 353 2267 388 2301
rect 422 2267 457 2301
rect 491 2267 526 2301
rect 560 2267 595 2301
rect 629 2267 664 2301
rect 698 2267 733 2301
rect 767 2267 802 2301
rect 836 2267 871 2301
rect 905 2267 940 2301
rect 974 2267 1009 2301
rect 1043 2267 1078 2301
rect 1112 2267 1146 2301
rect 1180 2267 1214 2301
rect 1248 2267 1282 2301
rect 1316 2267 1350 2301
rect 1384 2267 1418 2301
rect 1452 2267 1486 2301
rect 1520 2267 1554 2301
rect 1588 2267 1622 2301
rect 1656 2267 1690 2301
rect 1724 2267 1758 2301
rect 1792 2267 1826 2301
rect 1860 2267 1894 2301
rect 1928 2267 1962 2301
rect 1996 2267 2030 2301
rect 2064 2267 2098 2301
rect 2132 2267 2166 2301
rect 2200 2267 2234 2301
rect 2268 2267 2302 2301
rect 2336 2267 2370 2301
rect 2404 2267 2438 2301
rect 2472 2267 2506 2301
rect 2540 2267 2574 2301
rect 2608 2267 2642 2301
rect 2676 2267 2710 2301
rect 2744 2267 2778 2301
rect 2812 2267 2846 2301
rect 2880 2267 2914 2301
rect 2948 2267 2982 2301
rect 3016 2267 3050 2301
rect 3084 2267 3118 2301
rect 3152 2267 3186 2301
rect 3220 2267 3254 2301
rect 3288 2267 3322 2301
rect 3356 2267 3390 2301
rect 3424 2267 3458 2301
rect 3492 2267 3526 2301
rect 3560 2267 3594 2301
rect 3628 2267 3662 2301
rect 3696 2267 3730 2301
rect 3764 2267 3798 2301
rect 3832 2267 3866 2301
rect 3900 2267 3934 2301
rect 3968 2267 4002 2301
rect 4036 2267 4070 2301
rect 4104 2267 4138 2301
rect 4172 2267 4206 2301
rect 4240 2267 4274 2301
rect 4308 2267 4342 2301
rect 4376 2267 4410 2301
rect 4444 2267 4478 2301
rect 4512 2267 4546 2301
rect 4580 2267 4614 2301
rect 4648 2267 4682 2301
rect 4716 2267 4750 2301
rect 4784 2267 4818 2301
rect 4852 2267 4886 2301
rect 4920 2267 4954 2301
rect 4988 2267 5022 2301
rect 5056 2267 5090 2301
rect 5124 2267 5158 2301
rect 5192 2267 5226 2301
rect 5260 2267 5294 2301
rect 5328 2267 5362 2301
rect 5396 2267 5430 2301
rect 5464 2267 5498 2301
rect 5532 2267 5566 2301
rect 5600 2267 5634 2301
rect 5668 2267 5702 2301
rect 5736 2267 5770 2301
rect 5804 2267 5838 2301
rect 5872 2267 5906 2301
rect 5940 2267 5974 2301
rect 6008 2267 6042 2301
rect 6076 2277 6168 2301
rect 6076 2267 6134 2277
rect 88 2191 122 2267
rect 6134 2208 6168 2243
rect 88 2118 122 2157
rect 88 2045 122 2084
rect 88 1972 122 2011
rect 88 1899 122 1938
rect 88 1827 122 1865
rect 88 1755 122 1793
rect 88 1683 122 1721
rect 88 1611 122 1649
rect 88 1539 122 1577
rect 88 1467 122 1505
rect 88 1395 122 1433
rect 88 1323 122 1361
rect 88 1251 122 1289
rect 88 1193 122 1217
rect 6134 2139 6168 2174
rect 6134 2070 6168 2105
rect 6134 2001 6168 2036
rect 6134 1932 6168 1967
rect 6134 1863 6168 1898
rect 6134 1795 6168 1829
rect 6134 1727 6168 1761
rect 6134 1659 6168 1693
rect 6134 1591 6168 1625
rect 6134 1523 6168 1557
rect 6134 1455 6168 1489
rect 6134 1387 6168 1421
rect 6134 1319 6168 1353
rect 6134 1251 6168 1285
rect 1280 1039 1304 1073
rect 1338 1039 1373 1073
rect 1407 1039 1442 1073
rect 1476 1039 1511 1073
rect 1545 1039 1580 1073
rect 1614 1039 1649 1073
rect 1683 1039 1718 1073
rect 1752 1039 1787 1073
rect 1821 1039 1856 1073
rect 1890 1039 1925 1073
rect 1959 1039 1994 1073
rect 2028 1039 2063 1073
rect 2097 1039 2132 1073
rect 2166 1039 2201 1073
rect 2235 1039 2270 1073
rect 2304 1039 2339 1073
rect 2373 1039 2408 1073
rect 2442 1039 2477 1073
rect 2511 1039 2546 1073
rect 2580 1039 2615 1073
rect 2649 1039 2683 1073
rect 2717 1039 2751 1073
rect 2785 1039 2819 1073
rect 2853 1039 2877 1073
rect 3270 1039 3294 1073
rect 3328 1039 3363 1073
rect 3397 1039 3432 1073
rect 3466 1039 3501 1073
rect 3535 1039 3570 1073
rect 3604 1039 3639 1073
rect 3673 1039 3708 1073
rect 3742 1039 3777 1073
rect 3811 1039 3846 1073
rect 3880 1039 3914 1073
rect 3948 1039 3982 1073
rect 4016 1039 4050 1073
rect 4084 1039 4118 1073
rect 4152 1039 4186 1073
rect 4220 1039 4254 1073
rect 4288 1039 4322 1073
rect 4356 1039 4390 1073
rect 4424 1039 4458 1073
rect 4492 1039 4526 1073
rect 4560 1039 4584 1073
rect 6134 1073 6168 1217
rect 5663 1039 5687 1073
rect 5721 1039 5758 1073
rect 5792 1039 5829 1073
rect 5863 1039 5900 1073
rect 5934 1039 5970 1073
rect 6004 1039 6040 1073
rect 6074 1039 6110 1073
rect 6144 1039 6168 1073
<< psubdiffcont >>
rect 45 821 79 855
rect 45 751 79 785
rect 45 681 79 715
rect 45 611 79 645
rect 45 541 79 575
rect 45 472 79 506
rect 45 403 79 437
rect 45 334 79 368
rect 45 265 79 299
rect 5734 821 5768 855
rect 5734 747 5768 781
rect 5734 673 5768 707
rect 5734 599 5768 633
rect 5734 525 5768 559
rect 5734 451 5768 485
rect 5734 377 5768 411
rect 5734 303 5768 337
rect 69 171 103 205
rect 147 171 181 205
rect 225 171 259 205
rect 302 171 336 205
rect 379 171 413 205
rect 456 171 490 205
rect 533 171 567 205
rect 610 171 644 205
rect 2092 171 2126 205
rect 2162 171 2196 205
rect 2232 171 2266 205
rect 2302 171 2336 205
rect 2372 171 2406 205
rect 2442 171 2476 205
rect 2512 171 2546 205
rect 2582 171 2616 205
rect 2651 171 2685 205
rect 2720 171 2754 205
rect 2789 171 2823 205
rect 2858 171 2892 205
rect 2927 171 2961 205
rect 2996 171 3030 205
rect 3065 171 3099 205
rect 3134 171 3168 205
rect 3203 171 3237 205
rect 3272 171 3306 205
rect 3341 171 3375 205
rect 3410 171 3444 205
rect 3479 171 3513 205
rect 3548 171 3582 205
rect 3617 171 3651 205
rect 3686 171 3720 205
rect 3755 171 3789 205
rect 3824 171 3858 205
rect 3893 171 3927 205
rect 3962 171 3996 205
rect 4031 171 4065 205
rect 4827 171 4861 205
rect 4901 171 4935 205
rect 4975 171 5009 205
rect 5049 171 5083 205
rect 5123 171 5157 205
rect 5197 171 5231 205
rect 5271 171 5305 205
rect 5345 171 5379 205
rect 5418 171 5452 205
rect 5491 171 5525 205
rect 5564 171 5598 205
rect 5637 171 5671 205
rect 5710 171 5744 205
<< mvnsubdiffcont >>
rect 112 2267 146 2301
rect 181 2267 215 2301
rect 250 2267 284 2301
rect 319 2267 353 2301
rect 388 2267 422 2301
rect 457 2267 491 2301
rect 526 2267 560 2301
rect 595 2267 629 2301
rect 664 2267 698 2301
rect 733 2267 767 2301
rect 802 2267 836 2301
rect 871 2267 905 2301
rect 940 2267 974 2301
rect 1009 2267 1043 2301
rect 1078 2267 1112 2301
rect 1146 2267 1180 2301
rect 1214 2267 1248 2301
rect 1282 2267 1316 2301
rect 1350 2267 1384 2301
rect 1418 2267 1452 2301
rect 1486 2267 1520 2301
rect 1554 2267 1588 2301
rect 1622 2267 1656 2301
rect 1690 2267 1724 2301
rect 1758 2267 1792 2301
rect 1826 2267 1860 2301
rect 1894 2267 1928 2301
rect 1962 2267 1996 2301
rect 2030 2267 2064 2301
rect 2098 2267 2132 2301
rect 2166 2267 2200 2301
rect 2234 2267 2268 2301
rect 2302 2267 2336 2301
rect 2370 2267 2404 2301
rect 2438 2267 2472 2301
rect 2506 2267 2540 2301
rect 2574 2267 2608 2301
rect 2642 2267 2676 2301
rect 2710 2267 2744 2301
rect 2778 2267 2812 2301
rect 2846 2267 2880 2301
rect 2914 2267 2948 2301
rect 2982 2267 3016 2301
rect 3050 2267 3084 2301
rect 3118 2267 3152 2301
rect 3186 2267 3220 2301
rect 3254 2267 3288 2301
rect 3322 2267 3356 2301
rect 3390 2267 3424 2301
rect 3458 2267 3492 2301
rect 3526 2267 3560 2301
rect 3594 2267 3628 2301
rect 3662 2267 3696 2301
rect 3730 2267 3764 2301
rect 3798 2267 3832 2301
rect 3866 2267 3900 2301
rect 3934 2267 3968 2301
rect 4002 2267 4036 2301
rect 4070 2267 4104 2301
rect 4138 2267 4172 2301
rect 4206 2267 4240 2301
rect 4274 2267 4308 2301
rect 4342 2267 4376 2301
rect 4410 2267 4444 2301
rect 4478 2267 4512 2301
rect 4546 2267 4580 2301
rect 4614 2267 4648 2301
rect 4682 2267 4716 2301
rect 4750 2267 4784 2301
rect 4818 2267 4852 2301
rect 4886 2267 4920 2301
rect 4954 2267 4988 2301
rect 5022 2267 5056 2301
rect 5090 2267 5124 2301
rect 5158 2267 5192 2301
rect 5226 2267 5260 2301
rect 5294 2267 5328 2301
rect 5362 2267 5396 2301
rect 5430 2267 5464 2301
rect 5498 2267 5532 2301
rect 5566 2267 5600 2301
rect 5634 2267 5668 2301
rect 5702 2267 5736 2301
rect 5770 2267 5804 2301
rect 5838 2267 5872 2301
rect 5906 2267 5940 2301
rect 5974 2267 6008 2301
rect 6042 2267 6076 2301
rect 6134 2243 6168 2277
rect 88 2157 122 2191
rect 88 2084 122 2118
rect 88 2011 122 2045
rect 88 1938 122 1972
rect 88 1865 122 1899
rect 88 1793 122 1827
rect 88 1721 122 1755
rect 88 1649 122 1683
rect 88 1577 122 1611
rect 88 1505 122 1539
rect 88 1433 122 1467
rect 88 1361 122 1395
rect 88 1289 122 1323
rect 88 1217 122 1251
rect 6134 2174 6168 2208
rect 6134 2105 6168 2139
rect 6134 2036 6168 2070
rect 6134 1967 6168 2001
rect 6134 1898 6168 1932
rect 6134 1829 6168 1863
rect 6134 1761 6168 1795
rect 6134 1693 6168 1727
rect 6134 1625 6168 1659
rect 6134 1557 6168 1591
rect 6134 1489 6168 1523
rect 6134 1421 6168 1455
rect 6134 1353 6168 1387
rect 6134 1285 6168 1319
rect 6134 1217 6168 1251
rect 1304 1039 1338 1073
rect 1373 1039 1407 1073
rect 1442 1039 1476 1073
rect 1511 1039 1545 1073
rect 1580 1039 1614 1073
rect 1649 1039 1683 1073
rect 1718 1039 1752 1073
rect 1787 1039 1821 1073
rect 1856 1039 1890 1073
rect 1925 1039 1959 1073
rect 1994 1039 2028 1073
rect 2063 1039 2097 1073
rect 2132 1039 2166 1073
rect 2201 1039 2235 1073
rect 2270 1039 2304 1073
rect 2339 1039 2373 1073
rect 2408 1039 2442 1073
rect 2477 1039 2511 1073
rect 2546 1039 2580 1073
rect 2615 1039 2649 1073
rect 2683 1039 2717 1073
rect 2751 1039 2785 1073
rect 2819 1039 2853 1073
rect 3294 1039 3328 1073
rect 3363 1039 3397 1073
rect 3432 1039 3466 1073
rect 3501 1039 3535 1073
rect 3570 1039 3604 1073
rect 3639 1039 3673 1073
rect 3708 1039 3742 1073
rect 3777 1039 3811 1073
rect 3846 1039 3880 1073
rect 3914 1039 3948 1073
rect 3982 1039 4016 1073
rect 4050 1039 4084 1073
rect 4118 1039 4152 1073
rect 4186 1039 4220 1073
rect 4254 1039 4288 1073
rect 4322 1039 4356 1073
rect 4390 1039 4424 1073
rect 4458 1039 4492 1073
rect 4526 1039 4560 1073
rect 5687 1039 5721 1073
rect 5758 1039 5792 1073
rect 5829 1039 5863 1073
rect 5900 1039 5934 1073
rect 5970 1039 6004 1073
rect 6040 1039 6074 1073
rect 6110 1039 6144 1073
<< poly >>
rect 405 2193 505 2219
rect 691 2193 791 2219
rect 847 2193 947 2219
rect 1003 2193 1103 2219
rect 1159 2193 1259 2219
rect 1425 2193 1525 2219
rect 1581 2193 1681 2219
rect 1737 2193 1837 2219
rect 1893 2193 1993 2219
rect 2049 2193 2149 2219
rect 2205 2193 2305 2219
rect 2361 2193 2461 2219
rect 2517 2193 2617 2219
rect 2673 2193 2773 2219
rect 2829 2193 2929 2219
rect 2985 2193 3085 2219
rect 3141 2193 3241 2219
rect 3297 2193 3417 2219
rect 3473 2193 3593 2219
rect 3649 2193 3769 2219
rect 3825 2193 3945 2219
rect 4001 2193 4121 2219
rect 4177 2193 4297 2219
rect 4353 2193 4473 2219
rect 4529 2193 4649 2219
rect 4815 2193 4915 2219
rect 4971 2193 5071 2219
rect 5127 2193 5227 2219
rect 5283 2193 5383 2219
rect 5439 2193 5539 2219
rect 5595 2193 5695 2219
rect 5751 2193 5851 2219
rect 5907 2193 6007 2219
rect 405 1142 505 1193
rect 405 1108 436 1142
rect 470 1108 505 1142
rect 405 1074 505 1108
rect 405 1040 436 1074
rect 470 1040 505 1074
rect 405 1006 505 1040
rect 405 972 436 1006
rect 470 972 505 1006
rect 405 905 505 972
rect 691 1129 791 1193
rect 847 1167 947 1193
rect 691 1095 720 1129
rect 754 1095 791 1129
rect 691 1061 791 1095
rect 691 1027 720 1061
rect 754 1027 791 1061
rect 691 905 791 1027
rect 867 1129 947 1167
rect 867 1095 890 1129
rect 924 1095 947 1129
rect 867 1061 947 1095
rect 867 1027 890 1061
rect 924 1027 947 1061
rect 1003 1145 1103 1193
rect 1003 1111 1036 1145
rect 1070 1111 1103 1145
rect 1003 1077 1103 1111
rect 1003 1043 1036 1077
rect 1070 1043 1103 1077
rect 1003 1027 1103 1043
rect 1159 1145 1259 1193
rect 1159 1111 1175 1145
rect 1209 1111 1259 1145
rect 1159 1077 1259 1111
rect 1425 1167 1525 1193
rect 1581 1167 1681 1193
rect 1737 1167 1837 1193
rect 1893 1167 1993 1193
rect 2049 1167 2149 1193
rect 2205 1167 2305 1193
rect 1425 1145 2305 1167
rect 1425 1111 1483 1145
rect 1517 1111 1551 1145
rect 1585 1111 1619 1145
rect 1653 1111 1687 1145
rect 1721 1111 1755 1145
rect 1789 1111 1823 1145
rect 1857 1111 1891 1145
rect 1925 1111 1959 1145
rect 1993 1111 2027 1145
rect 2061 1111 2095 1145
rect 2129 1111 2163 1145
rect 2197 1111 2231 1145
rect 2265 1111 2305 1145
rect 1425 1095 2305 1111
rect 2361 1167 2461 1193
rect 2517 1167 2617 1193
rect 2673 1167 2773 1193
rect 2829 1167 2929 1193
rect 2985 1167 3085 1193
rect 3141 1167 3241 1193
rect 2361 1145 3241 1167
rect 2361 1111 2419 1145
rect 2453 1111 2487 1145
rect 2521 1111 2555 1145
rect 2589 1111 2623 1145
rect 2657 1111 2691 1145
rect 2725 1111 2759 1145
rect 2793 1111 2827 1145
rect 2861 1111 2895 1145
rect 2929 1111 2963 1145
rect 2997 1111 3031 1145
rect 3065 1111 3099 1145
rect 3133 1111 3167 1145
rect 3201 1111 3241 1145
rect 2361 1095 3241 1111
rect 3297 1167 3417 1193
rect 3473 1167 3593 1193
rect 3649 1167 3769 1193
rect 3825 1167 3945 1193
rect 4001 1167 4121 1193
rect 4177 1167 4297 1193
rect 4353 1167 4473 1193
rect 4529 1167 4649 1193
rect 4815 1167 4915 1193
rect 4971 1167 5071 1193
rect 5127 1167 5227 1193
rect 5283 1167 5383 1193
rect 5439 1167 5539 1193
rect 5595 1167 5695 1193
rect 5751 1167 5851 1193
rect 5907 1167 6007 1193
rect 3297 1145 4773 1167
rect 3297 1111 3335 1145
rect 3369 1111 3403 1145
rect 3437 1111 3471 1145
rect 3505 1111 3539 1145
rect 3573 1111 3607 1145
rect 3641 1111 3675 1145
rect 3709 1111 3743 1145
rect 3777 1111 3811 1145
rect 3845 1111 3879 1145
rect 3913 1111 3947 1145
rect 3981 1111 4015 1145
rect 4049 1111 4083 1145
rect 4117 1111 4151 1145
rect 4185 1111 4219 1145
rect 4253 1111 4287 1145
rect 4321 1111 4355 1145
rect 4389 1111 4423 1145
rect 4457 1111 4491 1145
rect 4525 1111 4559 1145
rect 4593 1111 4627 1145
rect 4661 1111 4695 1145
rect 4729 1111 4773 1145
rect 3297 1095 4773 1111
rect 4815 1145 5385 1167
rect 4815 1111 4835 1145
rect 4869 1111 4903 1145
rect 4937 1111 4971 1145
rect 5005 1111 5039 1145
rect 5073 1111 5107 1145
rect 5141 1111 5175 1145
rect 5209 1111 5243 1145
rect 5277 1111 5311 1145
rect 5345 1111 5385 1145
rect 4815 1095 5385 1111
rect 1159 1043 1175 1077
rect 1209 1043 1259 1077
rect 1159 1027 1259 1043
rect 2899 1057 3241 1095
rect 867 985 947 1027
rect 2899 1023 2919 1057
rect 2953 1023 2987 1057
rect 3021 1023 3055 1057
rect 3089 1023 3123 1057
rect 3157 1023 3191 1057
rect 3225 1023 3241 1057
rect 4607 1053 4773 1095
rect 867 969 1515 985
rect 2899 977 3241 1023
rect 4607 1029 4903 1053
rect 867 935 900 969
rect 934 935 968 969
rect 1002 935 1036 969
rect 1070 935 1104 969
rect 1138 935 1172 969
rect 1206 935 1240 969
rect 1274 935 1308 969
rect 1342 935 1376 969
rect 1410 935 1444 969
rect 1478 935 1515 969
rect 867 905 1515 935
rect 405 879 525 905
rect 691 879 811 905
rect 867 879 987 905
rect 1043 879 1163 905
rect 1219 879 1339 905
rect 1395 879 1515 905
rect 1681 961 1977 977
rect 1681 927 1717 961
rect 1751 927 1785 961
rect 1819 927 1853 961
rect 1887 927 1921 961
rect 1955 927 1977 961
rect 1681 905 1977 927
rect 1681 879 1801 905
rect 1857 879 1977 905
rect 2033 961 2329 977
rect 2033 927 2064 961
rect 2098 927 2132 961
rect 2166 927 2200 961
rect 2234 927 2268 961
rect 2302 927 2329 961
rect 2033 905 2329 927
rect 2033 879 2153 905
rect 2209 879 2329 905
rect 2495 961 3495 977
rect 2495 927 2545 961
rect 2579 927 2613 961
rect 2647 927 2681 961
rect 2715 927 2749 961
rect 2783 927 2817 961
rect 2851 927 2885 961
rect 2919 927 2953 961
rect 2987 927 3021 961
rect 3055 927 3089 961
rect 3123 927 3157 961
rect 3191 927 3225 961
rect 3259 927 3293 961
rect 3327 927 3361 961
rect 3395 927 3429 961
rect 3463 927 3495 961
rect 2495 905 3495 927
rect 2495 879 2615 905
rect 2671 879 2791 905
rect 2847 879 2967 905
rect 3023 879 3143 905
rect 3199 879 3319 905
rect 3375 879 3495 905
rect 3551 961 4551 977
rect 3551 927 3595 961
rect 3629 927 3663 961
rect 3697 927 3731 961
rect 3765 927 3799 961
rect 3833 927 3867 961
rect 3901 927 3935 961
rect 3969 927 4003 961
rect 4037 927 4071 961
rect 4105 927 4139 961
rect 4173 927 4207 961
rect 4241 927 4275 961
rect 4309 927 4343 961
rect 4377 927 4411 961
rect 4445 927 4479 961
rect 4513 927 4551 961
rect 3551 905 4551 927
rect 3551 879 3671 905
rect 3727 879 3847 905
rect 3903 879 4023 905
rect 4079 879 4199 905
rect 4255 879 4375 905
rect 4431 879 4551 905
rect 4607 927 4634 1029
rect 4872 927 4903 1029
rect 4607 905 4903 927
rect 4607 879 4727 905
rect 4783 879 4903 905
rect 4959 1029 5385 1095
rect 4959 927 4986 1029
rect 5224 1019 5385 1029
rect 5439 1145 6007 1167
rect 5439 1077 5471 1145
rect 5641 1111 5675 1145
rect 5709 1111 5743 1145
rect 5777 1111 5811 1145
rect 5845 1111 5879 1145
rect 5913 1111 5947 1145
rect 5981 1111 6007 1145
rect 5625 1095 6007 1111
rect 5439 1043 5455 1077
rect 5625 1043 5641 1095
rect 5224 927 5255 1019
rect 5439 977 5641 1043
rect 4959 905 5255 927
rect 4959 879 5079 905
rect 5135 879 5255 905
rect 5311 961 5641 977
rect 5311 927 5338 961
rect 5372 927 5406 961
rect 5440 927 5474 961
rect 5508 927 5542 961
rect 5576 927 5641 961
rect 5311 905 5641 927
rect 5311 879 5431 905
rect 5487 879 5607 905
rect 405 253 525 279
rect 691 253 811 279
rect 867 253 987 279
rect 1043 253 1163 279
rect 1219 253 1339 279
rect 1395 253 1515 279
rect 1681 253 1801 279
rect 1857 253 1977 279
rect 2033 253 2153 279
rect 2209 253 2329 279
rect 2495 253 2615 279
rect 2671 253 2791 279
rect 2847 253 2967 279
rect 3023 253 3143 279
rect 3199 253 3319 279
rect 3375 253 3495 279
rect 3551 253 3671 279
rect 3727 253 3847 279
rect 3903 253 4023 279
rect 4079 253 4199 279
rect 4255 253 4375 279
rect 4431 253 4551 279
rect 4607 253 4727 279
rect 4783 253 4903 279
rect 4959 253 5079 279
rect 5135 253 5255 279
rect 5311 253 5431 279
rect 5487 253 5607 279
<< polycont >>
rect 436 1108 470 1142
rect 436 1040 470 1074
rect 436 972 470 1006
rect 720 1095 754 1129
rect 720 1027 754 1061
rect 890 1095 924 1129
rect 890 1027 924 1061
rect 1036 1111 1070 1145
rect 1036 1043 1070 1077
rect 1175 1111 1209 1145
rect 1483 1111 1517 1145
rect 1551 1111 1585 1145
rect 1619 1111 1653 1145
rect 1687 1111 1721 1145
rect 1755 1111 1789 1145
rect 1823 1111 1857 1145
rect 1891 1111 1925 1145
rect 1959 1111 1993 1145
rect 2027 1111 2061 1145
rect 2095 1111 2129 1145
rect 2163 1111 2197 1145
rect 2231 1111 2265 1145
rect 2419 1111 2453 1145
rect 2487 1111 2521 1145
rect 2555 1111 2589 1145
rect 2623 1111 2657 1145
rect 2691 1111 2725 1145
rect 2759 1111 2793 1145
rect 2827 1111 2861 1145
rect 2895 1111 2929 1145
rect 2963 1111 2997 1145
rect 3031 1111 3065 1145
rect 3099 1111 3133 1145
rect 3167 1111 3201 1145
rect 3335 1111 3369 1145
rect 3403 1111 3437 1145
rect 3471 1111 3505 1145
rect 3539 1111 3573 1145
rect 3607 1111 3641 1145
rect 3675 1111 3709 1145
rect 3743 1111 3777 1145
rect 3811 1111 3845 1145
rect 3879 1111 3913 1145
rect 3947 1111 3981 1145
rect 4015 1111 4049 1145
rect 4083 1111 4117 1145
rect 4151 1111 4185 1145
rect 4219 1111 4253 1145
rect 4287 1111 4321 1145
rect 4355 1111 4389 1145
rect 4423 1111 4457 1145
rect 4491 1111 4525 1145
rect 4559 1111 4593 1145
rect 4627 1111 4661 1145
rect 4695 1111 4729 1145
rect 4835 1111 4869 1145
rect 4903 1111 4937 1145
rect 4971 1111 5005 1145
rect 5039 1111 5073 1145
rect 5107 1111 5141 1145
rect 5175 1111 5209 1145
rect 5243 1111 5277 1145
rect 5311 1111 5345 1145
rect 1175 1043 1209 1077
rect 2919 1023 2953 1057
rect 2987 1023 3021 1057
rect 3055 1023 3089 1057
rect 3123 1023 3157 1057
rect 3191 1023 3225 1057
rect 900 935 934 969
rect 968 935 1002 969
rect 1036 935 1070 969
rect 1104 935 1138 969
rect 1172 935 1206 969
rect 1240 935 1274 969
rect 1308 935 1342 969
rect 1376 935 1410 969
rect 1444 935 1478 969
rect 1717 927 1751 961
rect 1785 927 1819 961
rect 1853 927 1887 961
rect 1921 927 1955 961
rect 2064 927 2098 961
rect 2132 927 2166 961
rect 2200 927 2234 961
rect 2268 927 2302 961
rect 2545 927 2579 961
rect 2613 927 2647 961
rect 2681 927 2715 961
rect 2749 927 2783 961
rect 2817 927 2851 961
rect 2885 927 2919 961
rect 2953 927 2987 961
rect 3021 927 3055 961
rect 3089 927 3123 961
rect 3157 927 3191 961
rect 3225 927 3259 961
rect 3293 927 3327 961
rect 3361 927 3395 961
rect 3429 927 3463 961
rect 3595 927 3629 961
rect 3663 927 3697 961
rect 3731 927 3765 961
rect 3799 927 3833 961
rect 3867 927 3901 961
rect 3935 927 3969 961
rect 4003 927 4037 961
rect 4071 927 4105 961
rect 4139 927 4173 961
rect 4207 927 4241 961
rect 4275 927 4309 961
rect 4343 927 4377 961
rect 4411 927 4445 961
rect 4479 927 4513 961
rect 4634 927 4872 1029
rect 4986 927 5224 1029
rect 5471 1111 5641 1145
rect 5675 1111 5709 1145
rect 5743 1111 5777 1145
rect 5811 1111 5845 1145
rect 5879 1111 5913 1145
rect 5947 1111 5981 1145
rect 5471 1077 5625 1111
rect 5455 1043 5625 1077
rect 5338 927 5372 961
rect 5406 927 5440 961
rect 5474 927 5508 961
rect 5542 927 5576 961
<< locali >>
rect 88 2267 112 2301
rect 146 2267 181 2301
rect 215 2267 250 2301
rect 284 2267 319 2301
rect 353 2267 388 2301
rect 422 2267 457 2301
rect 491 2267 526 2301
rect 560 2267 595 2301
rect 629 2267 664 2301
rect 698 2267 733 2301
rect 767 2267 802 2301
rect 836 2267 871 2301
rect 905 2267 940 2301
rect 974 2267 1009 2301
rect 1043 2267 1078 2301
rect 1112 2267 1146 2301
rect 1180 2267 1214 2301
rect 1248 2267 1282 2301
rect 1316 2267 1350 2301
rect 1384 2267 1418 2301
rect 1452 2267 1486 2301
rect 1520 2267 1554 2301
rect 1588 2267 1622 2301
rect 1656 2267 1690 2301
rect 1724 2267 1758 2301
rect 1792 2267 1826 2301
rect 1860 2267 1894 2301
rect 1928 2267 1962 2301
rect 1996 2267 2030 2301
rect 2064 2267 2098 2301
rect 2132 2267 2166 2301
rect 2200 2267 2234 2301
rect 2268 2267 2302 2301
rect 2336 2267 2370 2301
rect 2404 2267 2438 2301
rect 2472 2267 2506 2301
rect 2540 2267 2574 2301
rect 2608 2267 2642 2301
rect 2676 2267 2710 2301
rect 2744 2267 2778 2301
rect 2812 2267 2846 2301
rect 2880 2267 2914 2301
rect 2948 2267 2982 2301
rect 3016 2267 3050 2301
rect 3084 2267 3118 2301
rect 3152 2267 3186 2301
rect 3220 2267 3254 2301
rect 3288 2267 3322 2301
rect 3356 2267 3390 2301
rect 3424 2267 3458 2301
rect 3492 2267 3526 2301
rect 3560 2267 3594 2301
rect 3628 2267 3662 2301
rect 3696 2267 3730 2301
rect 3764 2267 3798 2301
rect 3832 2267 3866 2301
rect 3900 2267 3934 2301
rect 3968 2267 4002 2301
rect 4036 2267 4070 2301
rect 4104 2267 4138 2301
rect 4172 2267 4206 2301
rect 4240 2267 4274 2301
rect 88 2223 122 2267
rect 88 2151 122 2157
rect 88 2079 122 2084
rect 88 1972 122 2011
rect 88 1899 122 1938
rect 88 1827 122 1865
rect 88 1755 122 1793
rect 88 1683 122 1721
rect 88 1611 122 1649
rect 88 1539 122 1577
rect 88 1467 122 1505
rect 88 1395 122 1433
rect 88 1323 122 1361
rect 88 1251 122 1289
rect 360 2223 394 2267
rect 802 2223 836 2267
rect 360 2181 394 2189
rect 360 2113 394 2117
rect 360 1977 394 2011
rect 360 1909 394 1943
rect 360 1841 394 1875
rect 360 1773 394 1807
rect 360 1705 394 1739
rect 360 1637 394 1671
rect 360 1569 394 1603
rect 360 1501 394 1535
rect 360 1433 394 1467
rect 360 1365 394 1399
rect 360 1297 394 1331
rect 360 1247 394 1263
rect 516 2181 570 2197
rect 550 2147 570 2181
rect 516 2113 570 2147
rect 550 2079 570 2113
rect 516 2045 570 2079
rect 550 2011 570 2045
rect 516 1977 570 2011
rect 550 1943 570 1977
rect 516 1909 570 1943
rect 550 1875 570 1909
rect 516 1841 570 1875
rect 550 1807 570 1841
rect 516 1773 570 1807
rect 550 1739 570 1773
rect 516 1705 570 1739
rect 550 1671 570 1705
rect 516 1637 570 1671
rect 550 1603 570 1637
rect 516 1569 570 1603
rect 550 1535 570 1569
rect 516 1501 570 1535
rect 550 1467 570 1501
rect 516 1433 570 1467
rect 550 1399 570 1433
rect 516 1365 570 1399
rect 550 1331 570 1365
rect 516 1297 570 1331
rect 550 1263 570 1297
rect 516 1228 570 1263
rect 88 1193 122 1217
rect 498 1194 536 1228
rect 436 1154 470 1158
rect 230 1120 268 1154
rect 302 1120 340 1154
rect 374 1120 412 1154
rect 446 1142 470 1154
rect 436 1074 470 1108
rect 436 1006 470 1040
rect 436 956 470 972
rect 45 855 79 879
rect 45 785 79 821
rect 45 734 79 751
rect 7 715 79 734
rect 7 681 45 715
rect 7 645 79 681
rect 7 611 45 645
rect 7 575 79 611
rect 7 541 45 575
rect 7 506 79 541
rect 7 484 45 506
rect 45 437 79 472
rect 45 368 79 403
rect 45 299 79 334
rect 360 761 394 767
rect 360 689 394 699
rect 360 597 394 631
rect 360 529 394 563
rect 360 461 394 495
rect 360 393 394 427
rect 360 325 394 359
rect 360 275 394 291
rect 516 801 570 1194
rect 516 767 536 801
rect 516 733 570 767
rect 516 699 536 733
rect 516 665 570 699
rect 516 631 536 665
rect 516 597 570 631
rect 516 563 536 597
rect 516 529 570 563
rect 516 495 536 529
rect 516 461 570 495
rect 516 427 536 461
rect 516 393 570 427
rect 516 359 536 393
rect 516 325 570 359
rect 516 291 536 325
rect 516 275 570 291
rect 622 2181 680 2197
rect 622 2147 646 2181
rect 622 2113 680 2147
rect 622 2079 646 2113
rect 622 2045 680 2079
rect 622 2011 646 2045
rect 622 1977 680 2011
rect 622 1943 646 1977
rect 622 1909 680 1943
rect 622 1875 646 1909
rect 622 1841 680 1875
rect 622 1807 646 1841
rect 622 1773 680 1807
rect 622 1739 646 1773
rect 622 1705 680 1739
rect 622 1671 646 1705
rect 622 1637 680 1671
rect 622 1603 646 1637
rect 622 1569 680 1603
rect 622 1535 646 1569
rect 622 1501 680 1535
rect 622 1467 646 1501
rect 622 1433 680 1467
rect 622 1399 646 1433
rect 622 1365 680 1399
rect 622 1331 646 1365
rect 622 1297 680 1331
rect 622 1263 646 1297
rect 622 1213 680 1263
rect 1114 2223 1148 2267
rect 802 2181 836 2189
rect 802 2113 836 2117
rect 802 1977 836 2011
rect 802 1909 836 1943
rect 802 1841 836 1875
rect 802 1773 836 1807
rect 802 1705 836 1739
rect 802 1637 836 1671
rect 802 1569 836 1603
rect 802 1501 836 1535
rect 802 1433 836 1467
rect 802 1365 836 1399
rect 802 1297 836 1331
rect 802 1247 836 1263
rect 958 2181 992 2197
rect 958 2113 992 2147
rect 958 2045 992 2079
rect 958 1977 992 2011
rect 958 1909 992 1943
rect 958 1841 992 1875
rect 958 1773 992 1807
rect 958 1705 992 1707
rect 958 1653 992 1671
rect 958 1569 992 1603
rect 958 1501 992 1532
rect 958 1433 992 1467
rect 958 1365 992 1399
rect 958 1297 992 1331
rect 958 1247 992 1263
rect 1380 2223 1414 2267
rect 1114 2181 1148 2189
rect 1114 2113 1148 2117
rect 1114 1977 1148 2011
rect 1114 1909 1148 1943
rect 1114 1841 1148 1875
rect 1114 1773 1148 1807
rect 1114 1705 1148 1739
rect 1114 1637 1148 1671
rect 1114 1569 1148 1603
rect 1114 1501 1148 1535
rect 1114 1433 1148 1467
rect 1114 1365 1148 1399
rect 1114 1297 1148 1331
rect 1114 1247 1148 1263
rect 1270 2181 1304 2197
rect 1270 2113 1304 2147
rect 1270 2045 1304 2079
rect 1270 1977 1304 2011
rect 1270 1909 1304 1943
rect 1270 1841 1304 1875
rect 1270 1773 1304 1807
rect 1270 1705 1304 1707
rect 1270 1653 1304 1671
rect 1270 1569 1304 1603
rect 1270 1501 1304 1532
rect 1270 1433 1304 1467
rect 1270 1365 1304 1399
rect 1270 1297 1304 1331
rect 622 1179 1070 1213
rect 622 913 680 1179
rect 1036 1145 1070 1179
rect 720 1129 754 1145
rect 720 1061 754 1095
rect 720 1011 754 1027
rect 890 1073 924 1095
rect 1036 1077 1070 1111
rect 1036 1027 1070 1039
rect 1175 1145 1209 1161
rect 1175 1077 1209 1111
rect 1270 1145 1304 1263
rect 1692 2223 1726 2267
rect 1380 2181 1414 2189
rect 1380 2113 1414 2117
rect 1380 1977 1414 2011
rect 1380 1909 1414 1943
rect 1380 1841 1414 1875
rect 1380 1773 1414 1807
rect 1380 1705 1414 1739
rect 1380 1637 1414 1671
rect 1380 1569 1414 1603
rect 1380 1501 1414 1535
rect 1380 1433 1414 1467
rect 1380 1365 1414 1399
rect 1380 1297 1414 1331
rect 1380 1247 1414 1263
rect 1536 2181 1570 2197
rect 1536 2113 1570 2147
rect 1536 2045 1570 2079
rect 2004 2223 2038 2267
rect 1692 2181 1726 2189
rect 1692 2113 1726 2117
rect 1536 1977 1570 2011
rect 1686 2011 1692 2033
rect 1848 2181 1882 2197
rect 1848 2113 1882 2147
rect 1848 2045 1882 2079
rect 1726 2011 1732 2033
rect 1686 2001 1732 2011
rect 1536 1940 1537 1943
rect 1536 1909 1571 1940
rect 1570 1897 1571 1909
rect 1536 1863 1537 1875
rect 1536 1841 1571 1863
rect 1570 1820 1571 1841
rect 1536 1786 1537 1807
rect 1536 1773 1571 1786
rect 1570 1743 1571 1773
rect 1536 1709 1537 1739
rect 1536 1705 1571 1709
rect 1570 1671 1571 1705
rect 1536 1666 1571 1671
rect 1536 1637 1537 1666
rect 1686 1943 1692 2001
rect 1726 1943 1732 2001
rect 1686 1925 1732 1943
rect 1686 1875 1692 1925
rect 1726 1875 1732 1925
rect 1686 1850 1732 1875
rect 1686 1807 1692 1850
rect 1726 1807 1732 1850
rect 1686 1775 1732 1807
rect 1686 1739 1692 1775
rect 1726 1739 1732 1775
rect 1686 1705 1732 1739
rect 1686 1666 1692 1705
rect 1726 1666 1732 1705
rect 1686 1637 1732 1666
rect 1686 1634 1692 1637
rect 1570 1603 1571 1632
rect 1536 1589 1571 1603
rect 1536 1569 1537 1589
rect 1726 1634 1732 1637
rect 2316 2223 2350 2267
rect 2004 2181 2038 2189
rect 2004 2113 2038 2117
rect 1848 1977 1882 2011
rect 1848 1909 1882 1940
rect 1848 1841 1882 1863
rect 1848 1773 1882 1786
rect 1848 1705 1882 1709
rect 1848 1666 1882 1671
rect 1692 1569 1726 1603
rect 1536 1501 1570 1535
rect 1536 1433 1570 1467
rect 1536 1365 1570 1399
rect 1536 1297 1570 1331
rect 1536 1247 1570 1263
rect 1692 1501 1726 1535
rect 1692 1433 1726 1467
rect 1692 1365 1726 1399
rect 1692 1297 1726 1331
rect 1692 1247 1726 1263
rect 1998 2011 2004 2033
rect 2160 2181 2194 2197
rect 2160 2113 2194 2147
rect 2160 2045 2194 2079
rect 2038 2011 2044 2033
rect 1998 2001 2044 2011
rect 1998 1943 2004 2001
rect 2038 1943 2044 2001
rect 1998 1925 2044 1943
rect 1998 1875 2004 1925
rect 2038 1875 2044 1925
rect 1998 1850 2044 1875
rect 1998 1807 2004 1850
rect 2038 1807 2044 1850
rect 1998 1775 2044 1807
rect 1998 1739 2004 1775
rect 2038 1739 2044 1775
rect 1998 1705 2044 1739
rect 1998 1666 2004 1705
rect 2038 1666 2044 1705
rect 1998 1637 2044 1666
rect 1998 1634 2004 1637
rect 1848 1589 1882 1603
rect 1848 1501 1882 1535
rect 1848 1433 1882 1467
rect 1848 1365 1882 1399
rect 1848 1297 1882 1331
rect 1848 1247 1882 1263
rect 2038 1634 2044 1637
rect 2628 2223 2662 2267
rect 2316 2181 2350 2189
rect 2316 2113 2350 2117
rect 2160 1977 2194 2011
rect 2160 1909 2194 1940
rect 2160 1841 2194 1863
rect 2160 1773 2194 1786
rect 2160 1705 2194 1709
rect 2160 1666 2194 1671
rect 2004 1569 2038 1603
rect 2004 1501 2038 1535
rect 2004 1433 2038 1467
rect 2004 1365 2038 1399
rect 2004 1297 2038 1331
rect 2004 1247 2038 1263
rect 2310 2011 2316 2033
rect 2472 2181 2506 2197
rect 2472 2113 2506 2147
rect 2472 2045 2506 2079
rect 2350 2011 2356 2033
rect 2310 2001 2356 2011
rect 2310 1943 2316 2001
rect 2350 1943 2356 2001
rect 2310 1925 2356 1943
rect 2310 1875 2316 1925
rect 2350 1875 2356 1925
rect 2310 1850 2356 1875
rect 2310 1807 2316 1850
rect 2350 1807 2356 1850
rect 2310 1775 2356 1807
rect 2310 1739 2316 1775
rect 2350 1739 2356 1775
rect 2310 1705 2356 1739
rect 2310 1666 2316 1705
rect 2350 1666 2356 1705
rect 2310 1637 2356 1666
rect 2310 1634 2316 1637
rect 2160 1589 2194 1603
rect 2160 1501 2194 1535
rect 2160 1433 2194 1467
rect 2160 1365 2194 1399
rect 2160 1297 2194 1331
rect 2160 1247 2194 1263
rect 2350 1634 2356 1637
rect 2940 2223 2974 2267
rect 2628 2181 2662 2189
rect 2628 2113 2662 2117
rect 2472 1977 2506 2011
rect 2472 1909 2506 1943
rect 2472 1841 2506 1875
rect 2472 1773 2506 1807
rect 2472 1705 2506 1739
rect 2472 1637 2506 1671
rect 2316 1569 2350 1603
rect 2316 1501 2350 1535
rect 2472 1569 2506 1603
rect 2622 2011 2628 2033
rect 2784 2181 2818 2197
rect 2784 2113 2818 2147
rect 2784 2045 2818 2079
rect 2662 2011 2668 2033
rect 2622 2001 2668 2011
rect 2622 1943 2628 2001
rect 2662 1943 2668 2001
rect 2622 1923 2668 1943
rect 2622 1875 2628 1923
rect 2662 1875 2668 1923
rect 2622 1845 2668 1875
rect 2622 1807 2628 1845
rect 2662 1807 2668 1845
rect 2622 1773 2668 1807
rect 2622 1733 2628 1773
rect 2662 1733 2668 1773
rect 2622 1705 2668 1733
rect 2622 1656 2628 1705
rect 2662 1656 2668 1705
rect 2622 1637 2668 1656
rect 2622 1579 2628 1637
rect 2662 1579 2668 1637
rect 2622 1569 2668 1579
rect 2622 1547 2628 1569
rect 2472 1501 2506 1535
rect 2316 1433 2350 1467
rect 2459 1467 2472 1473
rect 2662 1547 2668 1569
rect 3252 2223 3286 2267
rect 2940 2181 2974 2189
rect 2940 2113 2974 2117
rect 2784 1977 2818 2011
rect 2784 1939 2818 1943
rect 2784 1862 2818 1875
rect 2784 1785 2818 1807
rect 2784 1708 2818 1739
rect 2784 1637 2818 1671
rect 2934 2011 2940 2033
rect 3096 2181 3130 2197
rect 3096 2113 3130 2147
rect 3096 2045 3130 2079
rect 2974 2011 2980 2033
rect 2934 2001 2980 2011
rect 2934 1943 2940 2001
rect 2974 1943 2980 2001
rect 2934 1921 2980 1943
rect 2934 1875 2940 1921
rect 2974 1875 2980 1921
rect 2934 1842 2980 1875
rect 2934 1807 2940 1842
rect 2974 1807 2980 1842
rect 2934 1773 2980 1807
rect 2934 1729 2940 1773
rect 2974 1729 2980 1773
rect 2934 1705 2980 1729
rect 2934 1650 2940 1705
rect 2974 1650 2980 1705
rect 2934 1637 2980 1650
rect 2934 1618 2940 1637
rect 2784 1569 2818 1598
rect 2628 1501 2662 1535
rect 2506 1467 2519 1473
rect 2459 1439 2519 1467
rect 2316 1365 2350 1399
rect 2316 1297 2350 1331
rect 2316 1247 2350 1263
rect 2472 1433 2506 1439
rect 2472 1365 2506 1399
rect 2472 1297 2506 1331
rect 2472 1247 2506 1263
rect 2628 1433 2662 1467
rect 2628 1365 2662 1399
rect 2628 1297 2662 1331
rect 2628 1247 2662 1263
rect 2784 1501 2818 1522
rect 2784 1433 2818 1467
rect 2784 1365 2818 1399
rect 2784 1297 2818 1331
rect 2784 1247 2818 1263
rect 2974 1618 2980 1637
rect 3604 2223 3638 2267
rect 3252 2181 3286 2189
rect 3252 2113 3286 2117
rect 3096 1977 3130 2011
rect 3096 1939 3130 1943
rect 3246 2011 3252 2033
rect 3428 2181 3462 2197
rect 3428 2113 3462 2147
rect 3428 2045 3462 2079
rect 3286 2011 3292 2033
rect 3246 2001 3292 2011
rect 3246 1943 3252 2001
rect 3286 1943 3292 2001
rect 3096 1909 3097 1939
rect 3130 1875 3131 1905
rect 3096 1862 3131 1875
rect 3096 1841 3097 1862
rect 3130 1807 3131 1828
rect 3096 1785 3131 1807
rect 3096 1773 3097 1785
rect 3130 1739 3131 1751
rect 3096 1708 3131 1739
rect 3096 1705 3097 1708
rect 3130 1671 3131 1674
rect 3096 1637 3131 1671
rect 3130 1632 3131 1637
rect 2940 1569 2974 1603
rect 2940 1501 2974 1535
rect 2940 1433 2974 1467
rect 2940 1365 2974 1399
rect 2940 1297 2974 1331
rect 2940 1247 2974 1263
rect 3246 1921 3292 1943
rect 3246 1875 3252 1921
rect 3286 1875 3292 1921
rect 3246 1842 3292 1875
rect 3246 1807 3252 1842
rect 3286 1807 3292 1842
rect 3246 1773 3292 1807
rect 3246 1729 3252 1773
rect 3286 1729 3292 1773
rect 3246 1705 3292 1729
rect 3246 1650 3252 1705
rect 3286 1650 3292 1705
rect 3246 1637 3292 1650
rect 3246 1618 3252 1637
rect 3096 1598 3097 1603
rect 3096 1569 3131 1598
rect 3130 1556 3131 1569
rect 3096 1522 3097 1535
rect 3286 1618 3292 1637
rect 3956 2223 3990 2267
rect 3604 2181 3638 2189
rect 3604 2113 3638 2117
rect 3428 1977 3462 2011
rect 3428 1909 3462 1916
rect 3428 1873 3462 1875
rect 3428 1796 3462 1807
rect 3428 1719 3462 1739
rect 3428 1643 3462 1671
rect 3252 1569 3286 1603
rect 3096 1501 3130 1522
rect 3096 1433 3130 1467
rect 3096 1365 3130 1399
rect 3096 1297 3130 1331
rect 3096 1247 3130 1263
rect 3252 1501 3286 1535
rect 3252 1433 3286 1467
rect 3252 1365 3286 1399
rect 3252 1297 3286 1331
rect 3252 1247 3286 1263
rect 3598 2011 3604 2033
rect 3780 2181 3814 2197
rect 3780 2113 3814 2147
rect 3780 2045 3814 2079
rect 3638 2011 3644 2033
rect 3598 2001 3644 2011
rect 3598 1943 3604 2001
rect 3638 1943 3644 2001
rect 3598 1921 3644 1943
rect 3598 1875 3604 1921
rect 3638 1875 3644 1921
rect 3598 1842 3644 1875
rect 3598 1807 3604 1842
rect 3638 1807 3644 1842
rect 3598 1773 3644 1807
rect 3598 1729 3604 1773
rect 3638 1729 3644 1773
rect 3598 1705 3644 1729
rect 3598 1650 3604 1705
rect 3638 1650 3644 1705
rect 3598 1637 3644 1650
rect 3598 1618 3604 1637
rect 3428 1569 3462 1603
rect 3428 1501 3462 1533
rect 3428 1433 3462 1467
rect 3428 1365 3462 1399
rect 3428 1297 3462 1331
rect 3428 1247 3462 1263
rect 3638 1618 3644 1637
rect 4308 2223 4342 2301
rect 4376 2267 4410 2301
rect 4444 2267 4478 2301
rect 4512 2267 4546 2301
rect 4580 2267 4614 2301
rect 4648 2267 4682 2301
rect 4716 2267 4750 2301
rect 4784 2267 4818 2301
rect 4852 2267 4886 2301
rect 4920 2267 4954 2301
rect 4988 2267 5022 2301
rect 5056 2267 5090 2301
rect 5124 2267 5158 2301
rect 5192 2267 5226 2301
rect 5260 2267 5294 2301
rect 5328 2267 5362 2301
rect 5396 2267 5430 2301
rect 5464 2267 5498 2301
rect 5532 2267 5566 2301
rect 5600 2267 5634 2301
rect 5668 2267 5702 2301
rect 5736 2267 5770 2301
rect 5804 2267 5838 2301
rect 5872 2267 5906 2301
rect 5940 2267 5974 2301
rect 6008 2267 6042 2301
rect 6076 2277 6168 2301
rect 6076 2267 6134 2277
rect 3956 2181 3990 2189
rect 3956 2113 3990 2117
rect 3780 1977 3814 2011
rect 3780 1909 3814 1916
rect 3780 1873 3814 1875
rect 3780 1796 3814 1807
rect 3780 1719 3814 1739
rect 3780 1643 3814 1671
rect 3604 1569 3638 1603
rect 3604 1501 3638 1535
rect 3604 1433 3638 1467
rect 3604 1365 3638 1399
rect 3604 1297 3638 1331
rect 3604 1247 3638 1263
rect 3950 2011 3956 2033
rect 4132 2181 4166 2197
rect 4132 2113 4166 2147
rect 4132 2045 4166 2079
rect 3990 2011 3996 2033
rect 3950 2001 3996 2011
rect 3950 1943 3956 2001
rect 3990 1943 3996 2001
rect 3950 1921 3996 1943
rect 3950 1875 3956 1921
rect 3990 1875 3996 1921
rect 3950 1842 3996 1875
rect 3950 1807 3956 1842
rect 3990 1807 3996 1842
rect 3950 1773 3996 1807
rect 3950 1729 3956 1773
rect 3990 1729 3996 1773
rect 3950 1705 3996 1729
rect 3950 1650 3956 1705
rect 3990 1650 3996 1705
rect 3950 1637 3996 1650
rect 3950 1618 3956 1637
rect 3780 1569 3814 1603
rect 3780 1501 3814 1533
rect 3780 1433 3814 1467
rect 3780 1365 3814 1399
rect 3780 1297 3814 1331
rect 3780 1247 3814 1263
rect 3990 1618 3996 1637
rect 4660 2223 4694 2267
rect 4308 2181 4342 2189
rect 4308 2113 4342 2117
rect 4132 1977 4166 2011
rect 4132 1909 4166 1916
rect 4132 1873 4166 1875
rect 4132 1796 4166 1807
rect 4132 1719 4166 1739
rect 4132 1643 4166 1671
rect 3956 1569 3990 1603
rect 3956 1501 3990 1535
rect 3956 1433 3990 1467
rect 3956 1365 3990 1399
rect 3956 1297 3990 1331
rect 3956 1247 3990 1263
rect 4302 2011 4308 2033
rect 4484 2181 4518 2197
rect 4484 2113 4518 2147
rect 4484 2045 4518 2079
rect 4342 2011 4348 2033
rect 4302 2001 4348 2011
rect 4302 1943 4308 2001
rect 4342 1943 4348 2001
rect 4302 1921 4348 1943
rect 4302 1875 4308 1921
rect 4342 1875 4348 1921
rect 4302 1842 4348 1875
rect 4302 1807 4308 1842
rect 4342 1807 4348 1842
rect 4302 1773 4348 1807
rect 4302 1729 4308 1773
rect 4342 1729 4348 1773
rect 4302 1705 4348 1729
rect 4302 1650 4308 1705
rect 4342 1650 4348 1705
rect 4302 1637 4348 1650
rect 4302 1618 4308 1637
rect 4132 1569 4166 1603
rect 4132 1501 4166 1533
rect 4132 1433 4166 1467
rect 4132 1365 4166 1399
rect 4132 1297 4166 1331
rect 4132 1247 4166 1263
rect 4342 1618 4348 1637
rect 6134 2223 6168 2243
rect 4660 2181 4694 2189
rect 4660 2113 4694 2117
rect 4484 1977 4518 2011
rect 4484 1909 4518 1916
rect 4484 1873 4518 1875
rect 4484 1796 4518 1807
rect 4484 1719 4518 1739
rect 4484 1643 4518 1671
rect 4308 1569 4342 1603
rect 4308 1501 4342 1535
rect 4308 1433 4342 1467
rect 4308 1365 4342 1399
rect 4308 1297 4342 1331
rect 4308 1247 4342 1263
rect 4654 2011 4660 2033
rect 4770 2181 4804 2197
rect 4770 2113 4804 2147
rect 4770 2045 4804 2079
rect 4694 2011 4700 2033
rect 4654 2001 4700 2011
rect 4654 1943 4660 2001
rect 4694 1943 4700 2001
rect 4654 1921 4700 1943
rect 4654 1875 4660 1921
rect 4694 1875 4700 1921
rect 4654 1842 4700 1875
rect 4654 1807 4660 1842
rect 4694 1807 4700 1842
rect 4654 1773 4700 1807
rect 4654 1729 4660 1773
rect 4694 1729 4700 1773
rect 4654 1705 4700 1729
rect 4654 1650 4660 1705
rect 4694 1650 4700 1705
rect 4654 1637 4700 1650
rect 4654 1618 4660 1637
rect 4484 1569 4518 1603
rect 4484 1501 4518 1533
rect 4484 1433 4518 1467
rect 4484 1365 4518 1399
rect 4484 1297 4518 1331
rect 4484 1247 4518 1263
rect 4694 1618 4700 1637
rect 4770 1977 4804 2011
rect 4770 1909 4804 1939
rect 4770 1841 4804 1857
rect 4770 1773 4804 1775
rect 4770 1728 4804 1739
rect 4770 1647 4804 1671
rect 4660 1569 4694 1603
rect 4660 1501 4694 1535
rect 4660 1433 4694 1467
rect 4660 1365 4694 1399
rect 4660 1297 4694 1331
rect 4660 1247 4694 1263
rect 4770 1569 4804 1603
rect 4770 1501 4804 1535
rect 4770 1433 4804 1467
rect 4770 1365 4804 1399
rect 4770 1297 4804 1331
rect 4770 1247 4804 1263
rect 4926 2181 4960 2197
rect 4926 2113 4960 2147
rect 4926 2045 4960 2079
rect 4926 1977 4960 2011
rect 4926 1909 4960 1943
rect 4926 1869 4960 1875
rect 4926 1793 4960 1807
rect 4926 1717 4960 1739
rect 4926 1642 4960 1671
rect 4926 1569 4960 1603
rect 4926 1501 4960 1533
rect 4926 1433 4960 1467
rect 4926 1365 4960 1399
rect 4926 1297 4960 1331
rect 4926 1247 4960 1263
rect 5082 2181 5116 2197
rect 5082 2113 5116 2147
rect 5082 2045 5116 2079
rect 5082 1977 5116 2011
rect 5082 1909 5116 1939
rect 5082 1841 5116 1857
rect 5082 1773 5116 1775
rect 5082 1728 5116 1739
rect 5082 1647 5116 1671
rect 5082 1569 5116 1603
rect 5082 1501 5116 1535
rect 5082 1433 5116 1467
rect 5082 1365 5116 1399
rect 5082 1297 5116 1331
rect 5082 1247 5116 1263
rect 5238 2181 5272 2197
rect 5238 2113 5272 2147
rect 5238 2045 5272 2079
rect 5238 1977 5272 2011
rect 5238 1909 5272 1943
rect 5238 1869 5272 1875
rect 5394 2181 5428 2197
rect 5394 2113 5428 2147
rect 5394 2045 5428 2079
rect 5394 1977 5428 2011
rect 5394 1909 5428 1939
rect 5238 1841 5239 1869
rect 5272 1807 5273 1835
rect 5238 1783 5273 1807
rect 5238 1773 5239 1783
rect 5272 1739 5273 1749
rect 5238 1705 5273 1739
rect 5272 1698 5273 1705
rect 5238 1664 5239 1671
rect 5238 1637 5273 1664
rect 5272 1613 5273 1637
rect 5238 1579 5239 1603
rect 5238 1569 5273 1579
rect 5272 1535 5273 1569
rect 5238 1528 5273 1535
rect 5238 1501 5239 1528
rect 5272 1467 5273 1494
rect 5238 1443 5273 1467
rect 5238 1433 5239 1443
rect 5394 1841 5428 1863
rect 5394 1773 5428 1787
rect 5394 1705 5428 1711
rect 5394 1669 5428 1671
rect 5394 1593 5428 1603
rect 5394 1518 5428 1535
rect 5394 1443 5428 1467
rect 5238 1365 5272 1399
rect 5238 1297 5272 1331
rect 5238 1247 5272 1263
rect 5394 1365 5428 1399
rect 5394 1297 5428 1331
rect 5394 1247 5428 1263
rect 5550 2181 5584 2197
rect 5550 2113 5584 2147
rect 5550 2045 5584 2079
rect 5550 1977 5584 2011
rect 5550 1909 5584 1943
rect 5550 1841 5584 1853
rect 5550 1773 5584 1774
rect 5550 1729 5584 1739
rect 5550 1650 5584 1671
rect 5550 1571 5584 1603
rect 5550 1501 5584 1535
rect 5550 1433 5584 1459
rect 5550 1365 5584 1381
rect 5550 1297 5584 1303
rect 5550 1247 5584 1263
rect 5706 2181 5740 2197
rect 5706 2113 5740 2147
rect 5706 2045 5740 2079
rect 5706 1977 5740 2011
rect 5706 1909 5740 1939
rect 5706 1841 5740 1863
rect 5706 1773 5740 1787
rect 5706 1705 5740 1711
rect 5706 1669 5740 1671
rect 5706 1593 5740 1603
rect 5706 1518 5740 1535
rect 5706 1443 5740 1467
rect 5706 1365 5740 1399
rect 5706 1297 5740 1331
rect 5706 1247 5740 1263
rect 5862 2181 5896 2197
rect 5862 2113 5896 2147
rect 5862 2045 5896 2079
rect 5862 1977 5896 2011
rect 5862 1909 5896 1943
rect 5862 1841 5896 1853
rect 5862 1773 5896 1774
rect 5862 1729 5896 1739
rect 5862 1650 5896 1671
rect 5862 1572 5896 1603
rect 5862 1501 5896 1535
rect 5862 1433 5896 1460
rect 5862 1365 5896 1382
rect 5862 1297 5896 1304
rect 5862 1247 5896 1263
rect 6018 2181 6052 2197
rect 6018 2113 6052 2147
rect 6018 2045 6052 2079
rect 6018 1977 6052 2011
rect 6018 1909 6052 1939
rect 6018 1841 6052 1859
rect 6018 1773 6052 1780
rect 6018 1735 6052 1739
rect 6018 1656 6052 1671
rect 6018 1577 6052 1603
rect 6018 1501 6052 1535
rect 6018 1433 6052 1464
rect 6018 1365 6052 1385
rect 6018 1297 6052 1306
rect 6018 1247 6052 1263
rect 6168 2189 6206 2223
rect 6168 2174 6240 2189
rect 6134 2151 6240 2174
rect 6168 2137 6240 2151
rect 6168 2105 6206 2137
rect 6134 2103 6206 2105
rect 6134 2079 6240 2103
rect 6168 2051 6240 2079
rect 6168 2036 6206 2051
rect 6134 2017 6206 2036
rect 6134 2001 6240 2017
rect 6168 1967 6240 2001
rect 6134 1965 6240 1967
rect 6134 1932 6206 1965
rect 6168 1931 6206 1932
rect 6168 1898 6240 1931
rect 6134 1879 6240 1898
rect 6134 1863 6206 1879
rect 6168 1845 6206 1863
rect 6168 1829 6240 1845
rect 6134 1795 6240 1829
rect 6168 1773 6240 1795
rect 6134 1727 6168 1761
rect 6134 1659 6168 1692
rect 6134 1591 6168 1611
rect 6134 1523 6168 1529
rect 6134 1481 6168 1489
rect 6134 1399 6168 1421
rect 6134 1319 6168 1353
rect 6134 1251 6168 1283
rect 1270 1142 1483 1145
rect 1517 1142 1551 1145
rect 1585 1142 1619 1145
rect 1653 1142 1687 1145
rect 1721 1142 1755 1145
rect 1789 1142 1823 1145
rect 1857 1142 1891 1145
rect 1270 1108 1455 1142
rect 1517 1111 1527 1142
rect 1585 1111 1599 1142
rect 1653 1111 1671 1142
rect 1721 1111 1743 1142
rect 1789 1111 1815 1142
rect 1857 1111 1887 1142
rect 1925 1111 1959 1145
rect 1993 1111 2027 1145
rect 2061 1142 2095 1145
rect 2129 1142 2163 1145
rect 2197 1142 2231 1145
rect 2265 1142 2281 1145
rect 2403 1142 2419 1145
rect 2453 1142 2487 1145
rect 2521 1142 2555 1145
rect 2589 1142 2623 1145
rect 2657 1142 2691 1145
rect 2725 1142 2759 1145
rect 2793 1142 2827 1145
rect 2861 1142 2895 1145
rect 2065 1111 2095 1142
rect 2137 1111 2163 1142
rect 2209 1111 2231 1142
rect 1489 1108 1527 1111
rect 1561 1108 1599 1111
rect 1633 1108 1671 1111
rect 1705 1108 1743 1111
rect 1777 1108 1815 1111
rect 1849 1108 1887 1111
rect 1921 1108 1959 1111
rect 1993 1108 2031 1111
rect 2065 1108 2103 1111
rect 2137 1108 2175 1111
rect 2209 1108 2247 1111
rect 2453 1111 2459 1142
rect 2521 1111 2531 1142
rect 2589 1111 2603 1142
rect 2657 1111 2675 1142
rect 2725 1111 2747 1142
rect 2793 1111 2819 1142
rect 2861 1111 2891 1142
rect 2929 1111 2963 1145
rect 2997 1111 3031 1145
rect 3065 1142 3099 1145
rect 3133 1142 3167 1145
rect 3201 1142 3225 1145
rect 3069 1111 3099 1142
rect 3141 1111 3167 1142
rect 2421 1108 2459 1111
rect 2493 1108 2531 1111
rect 2565 1108 2603 1111
rect 2637 1108 2675 1111
rect 2709 1108 2747 1111
rect 2781 1108 2819 1111
rect 2853 1108 2891 1111
rect 2925 1108 2963 1111
rect 2997 1108 3035 1111
rect 3069 1108 3107 1111
rect 3141 1108 3179 1111
rect 3213 1108 3225 1142
rect 3319 1111 3335 1145
rect 3369 1142 3403 1145
rect 3437 1142 3471 1145
rect 3505 1142 3539 1145
rect 3573 1142 3607 1145
rect 3641 1142 3675 1145
rect 3384 1111 3403 1142
rect 3456 1111 3471 1142
rect 3528 1111 3539 1142
rect 3600 1111 3607 1142
rect 3672 1111 3675 1142
rect 3709 1142 3743 1145
rect 3777 1142 3811 1145
rect 3845 1142 3879 1145
rect 3913 1142 3947 1145
rect 3981 1142 4015 1145
rect 4049 1142 4083 1145
rect 4117 1142 4151 1145
rect 4185 1142 4219 1145
rect 4253 1142 4287 1145
rect 3709 1111 3710 1142
rect 3777 1111 3782 1142
rect 3845 1111 3854 1142
rect 3913 1111 3926 1142
rect 3981 1111 3998 1142
rect 4049 1111 4070 1142
rect 4117 1111 4142 1142
rect 4185 1111 4214 1142
rect 4253 1111 4286 1142
rect 4321 1111 4355 1145
rect 4389 1142 4423 1145
rect 4457 1142 4491 1145
rect 4525 1142 4559 1145
rect 4593 1142 4627 1145
rect 4661 1142 4695 1145
rect 4729 1142 4745 1145
rect 4819 1142 4835 1145
rect 4392 1111 4423 1142
rect 4464 1111 4491 1142
rect 4536 1111 4559 1142
rect 4608 1111 4627 1142
rect 4680 1111 4695 1142
rect 4819 1111 4831 1142
rect 4869 1111 4903 1145
rect 4937 1111 4971 1145
rect 5005 1142 5039 1145
rect 5073 1142 5107 1145
rect 5141 1142 5175 1145
rect 5209 1142 5243 1145
rect 5277 1142 5311 1145
rect 5345 1142 5361 1145
rect 5009 1111 5039 1142
rect 5081 1111 5107 1142
rect 5153 1111 5175 1142
rect 5225 1111 5243 1142
rect 5297 1111 5311 1142
rect 3384 1108 3422 1111
rect 3456 1108 3494 1111
rect 3528 1108 3566 1111
rect 3600 1108 3638 1111
rect 3672 1108 3710 1111
rect 3744 1108 3782 1111
rect 3816 1108 3854 1111
rect 3888 1108 3926 1111
rect 3960 1108 3998 1111
rect 4032 1108 4070 1111
rect 4104 1108 4142 1111
rect 4176 1108 4214 1111
rect 4248 1108 4286 1111
rect 4320 1108 4358 1111
rect 4392 1108 4430 1111
rect 4464 1108 4502 1111
rect 4536 1108 4574 1111
rect 4608 1108 4646 1111
rect 4680 1108 4718 1111
rect 4752 1108 4759 1111
rect 4865 1108 4903 1111
rect 4937 1108 4975 1111
rect 5009 1108 5047 1111
rect 5081 1108 5119 1111
rect 5153 1108 5191 1111
rect 5225 1108 5263 1111
rect 5297 1108 5335 1111
rect 1280 1062 1304 1073
rect 1338 1062 1373 1073
rect 1407 1062 1442 1073
rect 1476 1062 1511 1073
rect 1545 1062 1580 1073
rect 1280 1039 1289 1062
rect 1338 1039 1361 1062
rect 1407 1039 1433 1062
rect 1476 1039 1505 1062
rect 1545 1039 1577 1062
rect 1614 1039 1649 1073
rect 1683 1039 1718 1073
rect 1752 1062 1787 1073
rect 1821 1062 1856 1073
rect 1890 1062 1925 1073
rect 1959 1062 1994 1073
rect 2028 1062 2063 1073
rect 2097 1062 2132 1073
rect 2166 1062 2201 1073
rect 2235 1062 2270 1073
rect 2304 1062 2339 1073
rect 2373 1062 2408 1073
rect 2442 1062 2477 1073
rect 1755 1039 1787 1062
rect 1827 1039 1856 1062
rect 1899 1039 1925 1062
rect 1971 1039 1994 1062
rect 2043 1039 2063 1062
rect 2115 1039 2132 1062
rect 2187 1039 2201 1062
rect 2259 1039 2270 1062
rect 2331 1039 2339 1062
rect 2403 1039 2408 1062
rect 2475 1039 2477 1062
rect 2511 1062 2546 1073
rect 2580 1062 2615 1073
rect 2649 1062 2683 1073
rect 2717 1062 2751 1073
rect 2785 1062 2819 1073
rect 2511 1039 2513 1062
rect 2580 1039 2585 1062
rect 2649 1039 2657 1062
rect 2717 1039 2729 1062
rect 2785 1039 2801 1062
rect 2853 1039 2877 1073
rect 2919 1057 3225 1108
rect 1175 1027 1209 1039
rect 1323 1028 1361 1039
rect 1395 1028 1433 1039
rect 1467 1028 1505 1039
rect 1539 1028 1577 1039
rect 1611 1028 1649 1039
rect 1683 1028 1721 1039
rect 1755 1028 1793 1039
rect 1827 1028 1865 1039
rect 1899 1028 1937 1039
rect 1971 1028 2009 1039
rect 2043 1028 2081 1039
rect 2115 1028 2153 1039
rect 2187 1028 2225 1039
rect 2259 1028 2297 1039
rect 2331 1028 2369 1039
rect 2403 1028 2441 1039
rect 2475 1028 2513 1039
rect 2547 1028 2585 1039
rect 2619 1028 2657 1039
rect 2691 1028 2729 1039
rect 2763 1028 2801 1039
rect 890 969 924 1027
rect 2953 1023 2987 1057
rect 3021 1023 3055 1057
rect 3089 1023 3123 1057
rect 3157 1023 3191 1057
rect 3270 1039 3294 1073
rect 3328 1062 3363 1073
rect 3397 1062 3432 1073
rect 3466 1062 3501 1073
rect 3535 1062 3570 1073
rect 3604 1062 3639 1073
rect 3673 1062 3708 1073
rect 3742 1062 3777 1073
rect 3811 1062 3846 1073
rect 3880 1062 3914 1073
rect 3948 1062 3982 1073
rect 3332 1039 3363 1062
rect 3404 1039 3432 1062
rect 3476 1039 3501 1062
rect 3548 1039 3570 1062
rect 3620 1039 3639 1062
rect 3692 1039 3708 1062
rect 3764 1039 3777 1062
rect 3836 1039 3846 1062
rect 3908 1039 3914 1062
rect 3980 1039 3982 1062
rect 4016 1062 4050 1073
rect 4084 1062 4118 1073
rect 4152 1062 4186 1073
rect 4220 1062 4254 1073
rect 4288 1062 4322 1073
rect 4356 1062 4390 1073
rect 4424 1062 4458 1073
rect 4492 1062 4526 1073
rect 4016 1039 4018 1062
rect 4084 1039 4090 1062
rect 4152 1039 4162 1062
rect 4220 1039 4234 1062
rect 4288 1039 4306 1062
rect 4356 1039 4378 1062
rect 4424 1039 4450 1062
rect 4492 1039 4522 1062
rect 4560 1039 4584 1073
rect 3332 1028 3370 1039
rect 3404 1028 3442 1039
rect 3476 1028 3514 1039
rect 3548 1028 3586 1039
rect 3620 1028 3658 1039
rect 3692 1028 3730 1039
rect 3764 1028 3802 1039
rect 3836 1028 3874 1039
rect 3908 1028 3946 1039
rect 3980 1028 4018 1039
rect 4052 1028 4090 1039
rect 4124 1028 4162 1039
rect 4196 1028 4234 1039
rect 4268 1028 4306 1039
rect 4340 1028 4378 1039
rect 4412 1028 4450 1039
rect 4484 1028 4522 1039
rect 4618 1029 4759 1108
rect 4970 1029 5240 1108
rect 884 935 900 969
rect 934 935 968 969
rect 1002 935 1036 969
rect 1070 935 1104 969
rect 1138 935 1172 969
rect 1206 935 1240 969
rect 1274 935 1308 969
rect 1342 935 1376 969
rect 1410 935 1444 969
rect 1478 935 1494 969
rect 1701 954 1705 988
rect 1739 961 1777 988
rect 1811 961 1849 988
rect 1883 961 1921 988
rect 1751 954 1777 961
rect 1819 954 1849 961
rect 1701 927 1717 954
rect 1751 927 1785 954
rect 1819 927 1853 954
rect 1887 927 1921 961
rect 1955 927 1971 988
rect 2919 961 3225 1023
rect 2048 927 2064 961
rect 2098 927 2132 961
rect 2166 927 2200 961
rect 2234 927 2268 961
rect 2302 927 2318 961
rect 2529 927 2545 961
rect 2579 927 2613 961
rect 2647 927 2681 961
rect 2715 927 2749 961
rect 2783 927 2817 961
rect 2851 927 2885 961
rect 2919 927 2953 961
rect 2987 927 3021 961
rect 3055 927 3089 961
rect 3123 927 3157 961
rect 3191 927 3225 961
rect 3259 927 3293 961
rect 3327 927 3361 961
rect 3395 927 3429 961
rect 3463 927 3479 961
rect 3629 927 3635 961
rect 3697 927 3707 961
rect 3765 927 3779 961
rect 3833 927 3851 961
rect 3901 927 3923 961
rect 3969 927 3995 961
rect 4037 927 4067 961
rect 4105 927 4139 961
rect 4173 927 4207 961
rect 4245 927 4275 961
rect 4317 927 4343 961
rect 4377 927 4411 961
rect 4445 927 4479 961
rect 4513 927 4529 961
rect 4618 927 4634 1029
rect 4872 927 4888 1029
rect 4970 961 4986 1029
rect 5224 961 5240 1029
rect 5455 1077 5471 1145
rect 5641 1111 5675 1145
rect 5709 1111 5743 1145
rect 5777 1111 5811 1145
rect 5845 1111 5879 1145
rect 5913 1111 5947 1145
rect 5981 1111 5997 1145
rect 6134 1073 6168 1201
rect 5455 961 5625 1043
rect 5663 1062 5687 1073
rect 5721 1062 5758 1073
rect 5792 1062 5829 1073
rect 5863 1062 5900 1073
rect 5934 1062 5970 1073
rect 5721 1039 5735 1062
rect 5792 1039 5807 1062
rect 5863 1039 5879 1062
rect 5934 1039 5951 1062
rect 6004 1039 6040 1073
rect 6074 1039 6110 1073
rect 6144 1039 6168 1073
rect 5697 1028 5735 1039
rect 5769 1028 5807 1039
rect 5841 1028 5879 1039
rect 5913 1028 5951 1039
rect 4970 927 4978 961
rect 5228 927 5240 961
rect 5322 927 5338 961
rect 5372 927 5406 961
rect 5440 927 5474 961
rect 5508 927 5542 961
rect 5576 927 5625 961
rect 2048 913 2318 927
rect 656 879 694 913
rect 2082 879 2120 913
rect 2154 879 2192 913
rect 2226 879 2264 913
rect 2298 879 2318 913
rect 622 801 680 879
rect 5734 855 5768 879
rect 622 767 646 801
rect 622 733 680 767
rect 622 699 646 733
rect 622 665 680 699
rect 622 631 646 665
rect 822 761 856 767
rect 822 689 856 699
rect 622 597 680 631
rect 622 575 646 597
rect 622 541 634 575
rect 668 541 680 563
rect 622 529 680 541
rect 622 495 646 529
rect 622 461 634 495
rect 668 461 680 495
rect 622 427 646 461
rect 622 416 680 427
rect 622 382 634 416
rect 668 393 680 416
rect 622 359 646 382
rect 816 631 822 643
rect 998 801 1032 817
rect 998 733 1032 767
rect 998 665 1032 699
rect 856 631 862 643
rect 816 611 862 631
rect 816 563 822 611
rect 856 563 862 611
rect 816 529 862 563
rect 816 494 822 529
rect 856 494 862 529
rect 816 461 862 494
rect 816 412 822 461
rect 856 412 862 461
rect 816 393 862 412
rect 816 380 822 393
rect 622 337 680 359
rect 622 303 634 337
rect 668 325 680 337
rect 622 291 646 303
rect 622 275 680 291
rect 856 380 862 393
rect 1174 761 1208 767
rect 1174 689 1208 699
rect 998 597 1032 631
rect 998 529 1032 541
rect 998 416 1032 427
rect 822 325 856 359
rect 822 275 856 291
rect 1168 631 1174 643
rect 1350 801 1384 817
rect 1350 733 1384 767
rect 1350 665 1384 699
rect 1208 631 1214 643
rect 1168 611 1214 631
rect 1168 563 1174 611
rect 1208 563 1214 611
rect 1168 529 1214 563
rect 1168 494 1174 529
rect 1208 494 1214 529
rect 1168 461 1214 494
rect 1168 412 1174 461
rect 1208 412 1214 461
rect 1168 393 1214 412
rect 1168 380 1174 393
rect 998 337 1032 359
rect 998 275 1032 291
rect 1208 380 1214 393
rect 1526 761 1560 767
rect 1526 689 1560 699
rect 1350 597 1384 631
rect 1350 529 1384 541
rect 1350 416 1384 427
rect 1174 325 1208 359
rect 1174 275 1208 291
rect 1520 631 1526 643
rect 1636 801 1670 817
rect 1636 733 1670 767
rect 1636 665 1670 699
rect 1560 631 1566 643
rect 1520 611 1566 631
rect 1520 563 1526 611
rect 1560 563 1566 611
rect 1520 529 1566 563
rect 1520 494 1526 529
rect 1560 494 1566 529
rect 1520 461 1566 494
rect 1520 412 1526 461
rect 1560 412 1566 461
rect 1520 393 1566 412
rect 1520 380 1526 393
rect 1350 337 1384 359
rect 1350 275 1384 291
rect 1560 380 1566 393
rect 1636 597 1670 631
rect 1636 529 1670 562
rect 1636 461 1670 470
rect 1636 413 1670 427
rect 1526 325 1560 359
rect 1526 275 1560 291
rect 1636 325 1670 359
rect 1636 275 1670 291
rect 1812 801 1846 817
rect 1812 733 1846 767
rect 1812 665 1846 699
rect 1812 597 1846 631
rect 1812 529 1846 563
rect 1812 461 1846 482
rect 1812 426 1846 427
rect 1812 337 1846 359
rect 1812 275 1846 291
rect 1988 801 2022 817
rect 1988 733 2022 767
rect 1988 665 2022 699
rect 1988 597 2022 631
rect 1988 529 2022 562
rect 1988 461 2022 475
rect 1988 423 2022 427
rect 1988 337 2022 359
rect 1988 275 2022 291
rect 2164 801 2198 817
rect 2164 733 2198 767
rect 2164 665 2198 699
rect 2164 597 2198 631
rect 2164 529 2198 563
rect 2164 461 2198 482
rect 2164 426 2198 427
rect 2164 337 2198 359
rect 2164 275 2198 291
rect 2340 801 2374 817
rect 2340 733 2374 767
rect 2340 665 2374 699
rect 2450 761 2484 767
rect 2450 689 2484 699
rect 2340 597 2374 631
rect 2340 529 2374 562
rect 2340 461 2374 475
rect 2340 423 2374 427
rect 2340 337 2374 359
rect 2444 631 2450 643
rect 2626 801 2660 817
rect 2626 733 2660 767
rect 2626 665 2660 699
rect 2484 631 2490 643
rect 2444 611 2490 631
rect 2444 563 2450 611
rect 2484 563 2490 611
rect 2444 529 2490 563
rect 2444 492 2450 529
rect 2484 492 2490 529
rect 2444 461 2490 492
rect 2444 407 2450 461
rect 2484 407 2490 461
rect 2444 393 2490 407
rect 2444 359 2450 393
rect 2484 359 2490 393
rect 2444 357 2490 359
rect 2444 291 2450 357
rect 2484 291 2490 357
rect 2802 761 2836 767
rect 2802 689 2836 699
rect 2626 597 2660 631
rect 2626 529 2660 562
rect 2626 461 2660 475
rect 2626 423 2660 427
rect 2796 631 2802 643
rect 2978 801 3012 817
rect 2978 733 3012 767
rect 2978 665 3012 699
rect 2836 631 2842 643
rect 2796 611 2842 631
rect 2796 563 2802 611
rect 2836 563 2842 611
rect 2796 529 2842 563
rect 2796 494 2802 529
rect 2836 494 2842 529
rect 2796 461 2842 494
rect 2796 411 2802 461
rect 2836 411 2842 461
rect 2796 393 2842 411
rect 2796 379 2802 393
rect 2626 337 2660 359
rect 2340 275 2374 291
rect 2450 275 2484 291
rect 2626 275 2660 291
rect 2836 379 2842 393
rect 3154 761 3188 767
rect 3154 689 3188 699
rect 2978 597 3012 631
rect 2978 529 3012 562
rect 2978 461 3012 475
rect 2978 423 3012 427
rect 2802 325 2836 359
rect 2802 275 2836 291
rect 3148 631 3154 643
rect 3330 801 3364 817
rect 3330 733 3364 767
rect 3330 665 3364 699
rect 3188 631 3194 643
rect 3148 611 3194 631
rect 3148 563 3154 611
rect 3188 563 3194 611
rect 3148 529 3194 563
rect 3148 494 3154 529
rect 3188 494 3194 529
rect 3148 461 3194 494
rect 3148 411 3154 461
rect 3188 411 3194 461
rect 3148 393 3194 411
rect 3148 379 3154 393
rect 2978 337 3012 359
rect 2978 275 3012 291
rect 3188 379 3194 393
rect 3506 761 3540 767
rect 3506 689 3540 699
rect 3330 597 3364 631
rect 3330 529 3364 562
rect 3330 461 3364 475
rect 3330 423 3364 427
rect 3154 325 3188 359
rect 3154 275 3188 291
rect 3330 337 3364 359
rect 3330 275 3364 291
rect 3500 631 3506 643
rect 3682 801 3716 817
rect 3682 733 3716 767
rect 3682 665 3716 699
rect 3540 631 3546 643
rect 3500 611 3546 631
rect 3500 563 3506 611
rect 3540 563 3546 611
rect 3500 529 3546 563
rect 3500 487 3506 529
rect 3540 487 3546 529
rect 3500 461 3546 487
rect 3500 397 3506 461
rect 3540 397 3546 461
rect 3500 393 3546 397
rect 3500 359 3506 393
rect 3540 359 3546 393
rect 3500 341 3546 359
rect 3500 291 3506 341
rect 3540 291 3546 341
rect 3500 275 3546 291
rect 3858 761 3892 767
rect 3858 689 3892 699
rect 3682 597 3716 631
rect 3682 529 3716 562
rect 3682 461 3716 475
rect 3682 423 3716 427
rect 3852 631 3858 643
rect 4034 801 4068 817
rect 4034 733 4068 767
rect 4034 665 4068 699
rect 3892 631 3898 643
rect 3852 611 3898 631
rect 3852 563 3858 611
rect 3892 563 3898 611
rect 3852 529 3898 563
rect 3852 494 3858 529
rect 3892 494 3898 529
rect 3852 461 3898 494
rect 3852 411 3858 461
rect 3892 411 3898 461
rect 3852 393 3898 411
rect 3852 379 3858 393
rect 3682 337 3716 359
rect 3682 275 3716 291
rect 3892 379 3898 393
rect 4210 761 4244 767
rect 4210 689 4244 699
rect 4034 597 4068 631
rect 4034 529 4068 562
rect 4034 461 4068 475
rect 4034 423 4068 427
rect 3858 325 3892 359
rect 3858 275 3892 291
rect 4204 631 4210 643
rect 4386 801 4420 817
rect 4386 733 4420 767
rect 4386 665 4420 699
rect 4244 631 4250 643
rect 4204 611 4250 631
rect 4204 563 4210 611
rect 4244 563 4250 611
rect 4204 529 4250 563
rect 4204 494 4210 529
rect 4244 494 4250 529
rect 4204 461 4250 494
rect 4204 411 4210 461
rect 4244 411 4250 461
rect 4204 393 4250 411
rect 4204 379 4210 393
rect 4034 337 4068 359
rect 4034 275 4068 291
rect 4244 379 4250 393
rect 4386 597 4420 631
rect 4386 529 4420 562
rect 4386 461 4420 475
rect 4386 423 4420 427
rect 4210 325 4244 359
rect 4210 275 4244 291
rect 4386 337 4420 359
rect 4386 275 4420 291
rect 4562 761 4596 767
rect 4562 689 4596 699
rect 4562 597 4596 631
rect 4562 529 4596 563
rect 4562 461 4596 495
rect 4562 393 4596 427
rect 4562 325 4596 359
rect 4562 275 4596 291
rect 4738 801 4772 817
rect 4738 733 4772 767
rect 4738 665 4772 699
rect 4914 761 4948 767
rect 4914 689 4948 699
rect 4738 597 4772 631
rect 4738 529 4772 562
rect 4738 461 4772 475
rect 4738 423 4772 427
rect 4908 631 4914 643
rect 5090 801 5124 817
rect 5090 733 5124 767
rect 5090 665 5124 699
rect 4948 631 4954 643
rect 4908 611 4954 631
rect 4908 563 4914 611
rect 4948 563 4954 611
rect 4908 529 4954 563
rect 4908 494 4914 529
rect 4948 494 4954 529
rect 4908 461 4954 494
rect 4908 411 4914 461
rect 4948 411 4954 461
rect 4908 393 4954 411
rect 4908 379 4914 393
rect 4738 337 4772 359
rect 4738 275 4772 291
rect 4948 379 4954 393
rect 5266 761 5300 767
rect 5266 689 5300 699
rect 5090 597 5124 631
rect 5090 529 5124 562
rect 5090 461 5124 475
rect 5090 423 5124 427
rect 4914 325 4948 359
rect 4914 275 4948 291
rect 5260 631 5266 643
rect 5442 801 5476 817
rect 5442 733 5476 767
rect 5442 665 5476 699
rect 5300 631 5306 643
rect 5260 611 5306 631
rect 5260 563 5266 611
rect 5300 563 5306 611
rect 5260 529 5306 563
rect 5260 494 5266 529
rect 5300 494 5306 529
rect 5260 461 5306 494
rect 5260 411 5266 461
rect 5300 411 5306 461
rect 5260 393 5306 411
rect 5260 379 5266 393
rect 5090 337 5124 359
rect 5090 275 5124 291
rect 5300 379 5306 393
rect 5618 761 5652 767
rect 5618 689 5652 699
rect 5442 597 5476 631
rect 5442 529 5476 562
rect 5442 461 5476 475
rect 5442 423 5476 427
rect 5266 325 5300 359
rect 5266 275 5300 291
rect 5442 337 5476 359
rect 5442 275 5476 291
rect 5612 631 5618 643
rect 5734 781 5768 799
rect 5734 707 5768 727
rect 5652 631 5658 643
rect 5612 611 5658 631
rect 5612 563 5618 611
rect 5652 563 5658 611
rect 5612 529 5658 563
rect 5612 487 5618 529
rect 5652 487 5658 529
rect 5612 461 5658 487
rect 5612 397 5618 461
rect 5652 397 5658 461
rect 5612 393 5658 397
rect 5612 359 5618 393
rect 5652 359 5658 393
rect 5612 341 5658 359
rect 5612 291 5618 341
rect 5652 291 5658 341
rect 5612 275 5658 291
rect 5734 633 5768 655
rect 5734 559 5768 599
rect 5734 485 5768 525
rect 5734 411 5768 451
rect 5734 337 5768 377
rect 45 205 79 265
rect 5734 205 5768 303
rect 45 171 69 205
rect 103 171 147 205
rect 181 171 225 205
rect 259 171 302 205
rect 336 171 379 205
rect 413 171 456 205
rect 490 171 533 205
rect 567 171 610 205
rect 644 171 668 205
rect 2068 171 2092 205
rect 2126 171 2162 205
rect 2196 171 2232 205
rect 2266 171 2302 205
rect 2336 171 2372 205
rect 2406 171 2442 205
rect 2476 171 2512 205
rect 2546 171 2582 205
rect 2616 171 2651 205
rect 2685 171 2720 205
rect 2754 171 2789 205
rect 2823 171 2858 205
rect 2892 171 2927 205
rect 2961 171 2996 205
rect 3030 171 3065 205
rect 3099 171 3134 205
rect 3168 171 3203 205
rect 3237 171 3272 205
rect 3306 171 3341 205
rect 3375 171 3410 205
rect 3444 171 3479 205
rect 3513 171 3548 205
rect 3582 171 3617 205
rect 3651 171 3686 205
rect 3720 171 3755 205
rect 3789 171 3824 205
rect 3858 171 3893 205
rect 3927 171 3962 205
rect 3996 171 4031 205
rect 4065 171 4089 205
rect 4803 171 4827 205
rect 4861 171 4901 205
rect 4935 171 4975 205
rect 5009 171 5049 205
rect 5083 171 5123 205
rect 5157 171 5197 205
rect 5231 171 5271 205
rect 5305 171 5345 205
rect 5379 171 5418 205
rect 5452 171 5491 205
rect 5525 171 5564 205
rect 5598 171 5637 205
rect 5671 171 5710 205
rect 5744 171 5768 205
<< viali >>
rect 88 2191 122 2223
rect 88 2189 122 2191
rect 88 2118 122 2151
rect 88 2117 122 2118
rect 88 2045 122 2079
rect 360 2189 394 2223
rect 360 2147 394 2151
rect 360 2117 394 2147
rect 360 2045 394 2079
rect 464 1194 498 1228
rect 536 1194 570 1228
rect 196 1120 230 1154
rect 268 1120 302 1154
rect 340 1120 374 1154
rect 412 1142 446 1154
rect 412 1120 436 1142
rect 436 1120 446 1142
rect -99 484 7 734
rect 360 801 394 833
rect 360 799 394 801
rect 360 733 394 761
rect 360 727 394 733
rect 360 665 394 689
rect 360 655 394 665
rect 802 2189 836 2223
rect 802 2147 836 2151
rect 802 2117 836 2147
rect 802 2045 836 2079
rect 958 1739 992 1741
rect 958 1707 992 1739
rect 958 1637 992 1653
rect 958 1619 992 1637
rect 958 1535 992 1566
rect 958 1532 992 1535
rect 1114 2189 1148 2223
rect 1114 2147 1148 2151
rect 1114 2117 1148 2147
rect 1114 2045 1148 2079
rect 1270 1739 1304 1741
rect 1270 1707 1304 1739
rect 1270 1637 1304 1653
rect 1270 1619 1304 1637
rect 1270 1535 1304 1566
rect 1270 1532 1304 1535
rect 890 1129 924 1145
rect 890 1111 924 1129
rect 890 1061 924 1073
rect 890 1039 924 1061
rect 1036 1111 1070 1145
rect 1036 1043 1070 1073
rect 1036 1039 1070 1043
rect 1175 1111 1209 1145
rect 1380 2189 1414 2223
rect 1380 2147 1414 2151
rect 1380 2117 1414 2147
rect 1380 2045 1414 2079
rect 1692 2189 1726 2223
rect 1692 2147 1726 2151
rect 1692 2117 1726 2147
rect 1692 2045 1726 2079
rect 1537 1943 1570 1974
rect 1570 1943 1571 1974
rect 1537 1940 1571 1943
rect 1537 1875 1570 1897
rect 1570 1875 1571 1897
rect 1537 1863 1571 1875
rect 1537 1807 1570 1820
rect 1570 1807 1571 1820
rect 1537 1786 1571 1807
rect 1537 1739 1570 1743
rect 1570 1739 1571 1743
rect 1537 1709 1571 1739
rect 1537 1637 1571 1666
rect 1537 1632 1570 1637
rect 1570 1632 1571 1637
rect 1692 1977 1726 2001
rect 1692 1967 1726 1977
rect 1692 1909 1726 1925
rect 1692 1891 1726 1909
rect 1692 1841 1726 1850
rect 1692 1816 1726 1841
rect 1692 1773 1726 1775
rect 1692 1741 1726 1773
rect 1692 1671 1726 1700
rect 1692 1666 1726 1671
rect 1537 1569 1571 1589
rect 1537 1555 1570 1569
rect 1570 1555 1571 1569
rect 2004 2189 2038 2223
rect 2004 2147 2038 2151
rect 2004 2117 2038 2147
rect 2004 2045 2038 2079
rect 1848 1943 1882 1974
rect 1848 1940 1882 1943
rect 1848 1875 1882 1897
rect 1848 1863 1882 1875
rect 1848 1807 1882 1820
rect 1848 1786 1882 1807
rect 1848 1739 1882 1743
rect 1848 1709 1882 1739
rect 1848 1637 1882 1666
rect 1848 1632 1882 1637
rect 2004 1977 2038 2001
rect 2004 1967 2038 1977
rect 2004 1909 2038 1925
rect 2004 1891 2038 1909
rect 2004 1841 2038 1850
rect 2004 1816 2038 1841
rect 2004 1773 2038 1775
rect 2004 1741 2038 1773
rect 2004 1671 2038 1700
rect 2004 1666 2038 1671
rect 1848 1569 1882 1589
rect 1848 1555 1882 1569
rect 2316 2189 2350 2223
rect 2316 2147 2350 2151
rect 2316 2117 2350 2147
rect 2316 2045 2350 2079
rect 2160 1943 2194 1974
rect 2160 1940 2194 1943
rect 2160 1875 2194 1897
rect 2160 1863 2194 1875
rect 2160 1807 2194 1820
rect 2160 1786 2194 1807
rect 2160 1739 2194 1743
rect 2160 1709 2194 1739
rect 2160 1637 2194 1666
rect 2160 1632 2194 1637
rect 2316 1977 2350 2001
rect 2316 1967 2350 1977
rect 2316 1909 2350 1925
rect 2316 1891 2350 1909
rect 2316 1841 2350 1850
rect 2316 1816 2350 1841
rect 2316 1773 2350 1775
rect 2316 1741 2350 1773
rect 2316 1671 2350 1700
rect 2316 1666 2350 1671
rect 2160 1569 2194 1589
rect 2160 1555 2194 1569
rect 2628 2189 2662 2223
rect 2628 2147 2662 2151
rect 2628 2117 2662 2147
rect 2628 2045 2662 2079
rect 2628 1977 2662 2001
rect 2628 1967 2662 1977
rect 2628 1909 2662 1923
rect 2628 1889 2662 1909
rect 2628 1841 2662 1845
rect 2628 1811 2662 1841
rect 2628 1739 2662 1767
rect 2628 1733 2662 1739
rect 2628 1671 2662 1690
rect 2628 1656 2662 1671
rect 2628 1603 2662 1613
rect 2628 1579 2662 1603
rect 2425 1439 2459 1473
rect 2940 2189 2974 2223
rect 2940 2147 2974 2151
rect 2940 2117 2974 2147
rect 2940 2045 2974 2079
rect 2784 1909 2818 1939
rect 2784 1905 2818 1909
rect 2784 1841 2818 1862
rect 2784 1828 2818 1841
rect 2784 1773 2818 1785
rect 2784 1751 2818 1773
rect 2784 1705 2818 1708
rect 2784 1674 2818 1705
rect 2784 1603 2818 1632
rect 2940 1977 2974 2001
rect 2940 1967 2974 1977
rect 2940 1909 2974 1921
rect 2940 1887 2974 1909
rect 2940 1841 2974 1842
rect 2940 1808 2974 1841
rect 2940 1739 2974 1763
rect 2940 1729 2974 1739
rect 2940 1671 2974 1684
rect 2940 1650 2974 1671
rect 2784 1598 2818 1603
rect 2519 1439 2553 1473
rect 2784 1535 2818 1556
rect 2784 1522 2818 1535
rect 3252 2189 3286 2223
rect 3252 2147 3286 2151
rect 3252 2117 3286 2147
rect 3252 2045 3286 2079
rect 3252 1977 3286 2001
rect 3252 1967 3286 1977
rect 3097 1909 3131 1939
rect 3097 1905 3130 1909
rect 3130 1905 3131 1909
rect 3097 1841 3131 1862
rect 3097 1828 3130 1841
rect 3130 1828 3131 1841
rect 3097 1773 3131 1785
rect 3097 1751 3130 1773
rect 3130 1751 3131 1773
rect 3097 1705 3131 1708
rect 3097 1674 3130 1705
rect 3130 1674 3131 1705
rect 3097 1603 3130 1632
rect 3130 1603 3131 1632
rect 3252 1909 3286 1921
rect 3252 1887 3286 1909
rect 3252 1841 3286 1842
rect 3252 1808 3286 1841
rect 3252 1739 3286 1763
rect 3252 1729 3286 1739
rect 3252 1671 3286 1684
rect 3252 1650 3286 1671
rect 3097 1598 3131 1603
rect 3097 1535 3130 1556
rect 3130 1535 3131 1556
rect 3097 1522 3131 1535
rect 3604 2189 3638 2223
rect 3604 2147 3638 2151
rect 3604 2117 3638 2147
rect 3604 2045 3638 2079
rect 3428 1943 3462 1950
rect 3428 1916 3462 1943
rect 3428 1841 3462 1873
rect 3428 1839 3462 1841
rect 3428 1773 3462 1796
rect 3428 1762 3462 1773
rect 3428 1705 3462 1719
rect 3428 1685 3462 1705
rect 3428 1637 3462 1643
rect 3428 1609 3462 1637
rect 3604 1977 3638 2001
rect 3604 1967 3638 1977
rect 3604 1909 3638 1921
rect 3604 1887 3638 1909
rect 3604 1841 3638 1842
rect 3604 1808 3638 1841
rect 3604 1739 3638 1763
rect 3604 1729 3638 1739
rect 3604 1671 3638 1684
rect 3604 1650 3638 1671
rect 3428 1535 3462 1567
rect 3428 1533 3462 1535
rect 3956 2189 3990 2223
rect 3956 2147 3990 2151
rect 3956 2117 3990 2147
rect 3956 2045 3990 2079
rect 3780 1943 3814 1950
rect 3780 1916 3814 1943
rect 3780 1841 3814 1873
rect 3780 1839 3814 1841
rect 3780 1773 3814 1796
rect 3780 1762 3814 1773
rect 3780 1705 3814 1719
rect 3780 1685 3814 1705
rect 3780 1637 3814 1643
rect 3780 1609 3814 1637
rect 3956 1977 3990 2001
rect 3956 1967 3990 1977
rect 3956 1909 3990 1921
rect 3956 1887 3990 1909
rect 3956 1841 3990 1842
rect 3956 1808 3990 1841
rect 3956 1739 3990 1763
rect 3956 1729 3990 1739
rect 3956 1671 3990 1684
rect 3956 1650 3990 1671
rect 3780 1535 3814 1567
rect 3780 1533 3814 1535
rect 4308 2189 4342 2223
rect 4308 2147 4342 2151
rect 4308 2117 4342 2147
rect 4308 2045 4342 2079
rect 4132 1943 4166 1950
rect 4132 1916 4166 1943
rect 4132 1841 4166 1873
rect 4132 1839 4166 1841
rect 4132 1773 4166 1796
rect 4132 1762 4166 1773
rect 4132 1705 4166 1719
rect 4132 1685 4166 1705
rect 4132 1637 4166 1643
rect 4132 1609 4166 1637
rect 4308 1977 4342 2001
rect 4308 1967 4342 1977
rect 4308 1909 4342 1921
rect 4308 1887 4342 1909
rect 4308 1841 4342 1842
rect 4308 1808 4342 1841
rect 4308 1739 4342 1763
rect 4308 1729 4342 1739
rect 4308 1671 4342 1684
rect 4308 1650 4342 1671
rect 4132 1535 4166 1567
rect 4132 1533 4166 1535
rect 4660 2189 4694 2223
rect 6134 2208 6168 2223
rect 4660 2147 4694 2151
rect 4660 2117 4694 2147
rect 4660 2045 4694 2079
rect 4484 1943 4518 1950
rect 4484 1916 4518 1943
rect 4484 1841 4518 1873
rect 4484 1839 4518 1841
rect 4484 1773 4518 1796
rect 4484 1762 4518 1773
rect 4484 1705 4518 1719
rect 4484 1685 4518 1705
rect 4484 1637 4518 1643
rect 4484 1609 4518 1637
rect 4660 1977 4694 2001
rect 4660 1967 4694 1977
rect 4660 1909 4694 1921
rect 4660 1887 4694 1909
rect 4660 1841 4694 1842
rect 4660 1808 4694 1841
rect 4660 1739 4694 1763
rect 4660 1729 4694 1739
rect 4660 1671 4694 1684
rect 4660 1650 4694 1671
rect 4484 1535 4518 1567
rect 4484 1533 4518 1535
rect 4770 1943 4804 1973
rect 4770 1939 4804 1943
rect 4770 1875 4804 1891
rect 4770 1857 4804 1875
rect 4770 1807 4804 1809
rect 4770 1775 4804 1807
rect 4770 1705 4804 1728
rect 4770 1694 4804 1705
rect 4770 1637 4804 1647
rect 4770 1613 4804 1637
rect 4926 1841 4960 1869
rect 4926 1835 4960 1841
rect 4926 1773 4960 1793
rect 4926 1759 4960 1773
rect 4926 1705 4960 1717
rect 4926 1683 4960 1705
rect 4926 1637 4960 1642
rect 4926 1608 4960 1637
rect 4926 1535 4960 1567
rect 4926 1533 4960 1535
rect 5082 1943 5116 1973
rect 5082 1939 5116 1943
rect 5082 1875 5116 1891
rect 5082 1857 5116 1875
rect 5082 1807 5116 1809
rect 5082 1775 5116 1807
rect 5082 1705 5116 1728
rect 5082 1694 5116 1705
rect 5082 1637 5116 1647
rect 5082 1613 5116 1637
rect 5394 1943 5428 1973
rect 5394 1939 5428 1943
rect 5394 1875 5428 1897
rect 5239 1841 5273 1869
rect 5239 1835 5272 1841
rect 5272 1835 5273 1841
rect 5239 1773 5273 1783
rect 5239 1749 5272 1773
rect 5272 1749 5273 1773
rect 5239 1671 5272 1698
rect 5272 1671 5273 1698
rect 5239 1664 5273 1671
rect 5239 1603 5272 1613
rect 5272 1603 5273 1613
rect 5239 1579 5273 1603
rect 5239 1501 5273 1528
rect 5239 1494 5272 1501
rect 5272 1494 5273 1501
rect 5239 1433 5273 1443
rect 5239 1409 5272 1433
rect 5272 1409 5273 1433
rect 5394 1863 5428 1875
rect 5394 1807 5428 1821
rect 5394 1787 5428 1807
rect 5394 1739 5428 1745
rect 5394 1711 5428 1739
rect 5394 1637 5428 1669
rect 5394 1635 5428 1637
rect 5394 1569 5428 1593
rect 5394 1559 5428 1569
rect 5394 1501 5428 1518
rect 5394 1484 5428 1501
rect 5394 1433 5428 1443
rect 5394 1409 5428 1433
rect 5550 1875 5584 1887
rect 5550 1853 5584 1875
rect 5550 1807 5584 1808
rect 5550 1774 5584 1807
rect 5550 1705 5584 1729
rect 5550 1695 5584 1705
rect 5550 1637 5584 1650
rect 5550 1616 5584 1637
rect 5550 1569 5584 1571
rect 5550 1537 5584 1569
rect 5550 1467 5584 1493
rect 5550 1459 5584 1467
rect 5550 1399 5584 1415
rect 5550 1381 5584 1399
rect 5550 1331 5584 1337
rect 5550 1303 5584 1331
rect 5706 1943 5740 1973
rect 5706 1939 5740 1943
rect 5706 1875 5740 1897
rect 5706 1863 5740 1875
rect 5706 1807 5740 1821
rect 5706 1787 5740 1807
rect 5706 1739 5740 1745
rect 5706 1711 5740 1739
rect 5706 1637 5740 1669
rect 5706 1635 5740 1637
rect 5706 1569 5740 1593
rect 5706 1559 5740 1569
rect 5706 1501 5740 1518
rect 5706 1484 5740 1501
rect 5706 1433 5740 1443
rect 5706 1409 5740 1433
rect 5862 1875 5896 1887
rect 5862 1853 5896 1875
rect 5862 1807 5896 1808
rect 5862 1774 5896 1807
rect 5862 1705 5896 1729
rect 5862 1695 5896 1705
rect 5862 1637 5896 1650
rect 5862 1616 5896 1637
rect 5862 1569 5896 1572
rect 5862 1538 5896 1569
rect 5862 1467 5896 1494
rect 5862 1460 5896 1467
rect 5862 1399 5896 1416
rect 5862 1382 5896 1399
rect 5862 1331 5896 1338
rect 5862 1304 5896 1331
rect 6018 1943 6052 1973
rect 6018 1939 6052 1943
rect 6018 1875 6052 1893
rect 6018 1859 6052 1875
rect 6018 1807 6052 1814
rect 6018 1780 6052 1807
rect 6018 1705 6052 1735
rect 6018 1701 6052 1705
rect 6018 1637 6052 1656
rect 6018 1622 6052 1637
rect 6018 1569 6052 1577
rect 6018 1543 6052 1569
rect 6018 1467 6052 1498
rect 6018 1464 6052 1467
rect 6018 1399 6052 1419
rect 6018 1385 6052 1399
rect 6018 1331 6052 1340
rect 6018 1306 6052 1331
rect 6134 2189 6168 2208
rect 6206 2189 6240 2223
rect 6134 2139 6168 2151
rect 6134 2117 6168 2139
rect 6206 2103 6240 2137
rect 6134 2070 6168 2079
rect 6134 2045 6168 2070
rect 6206 2017 6240 2051
rect 6206 1931 6240 1965
rect 6206 1845 6240 1879
rect 6134 1693 6168 1726
rect 6134 1692 6168 1693
rect 6134 1625 6168 1645
rect 6134 1611 6168 1625
rect 6134 1557 6168 1563
rect 6134 1529 6168 1557
rect 6134 1455 6168 1481
rect 6134 1447 6168 1455
rect 6134 1387 6168 1399
rect 6134 1365 6168 1387
rect 6134 1285 6168 1317
rect 6134 1283 6168 1285
rect 6134 1217 6168 1235
rect 6134 1201 6168 1217
rect 1455 1111 1483 1142
rect 1483 1111 1489 1142
rect 1527 1111 1551 1142
rect 1551 1111 1561 1142
rect 1599 1111 1619 1142
rect 1619 1111 1633 1142
rect 1671 1111 1687 1142
rect 1687 1111 1705 1142
rect 1743 1111 1755 1142
rect 1755 1111 1777 1142
rect 1815 1111 1823 1142
rect 1823 1111 1849 1142
rect 1887 1111 1891 1142
rect 1891 1111 1921 1142
rect 1959 1111 1993 1142
rect 2031 1111 2061 1142
rect 2061 1111 2065 1142
rect 2103 1111 2129 1142
rect 2129 1111 2137 1142
rect 2175 1111 2197 1142
rect 2197 1111 2209 1142
rect 2247 1111 2265 1142
rect 2265 1111 2281 1142
rect 1455 1108 1489 1111
rect 1527 1108 1561 1111
rect 1599 1108 1633 1111
rect 1671 1108 1705 1111
rect 1743 1108 1777 1111
rect 1815 1108 1849 1111
rect 1887 1108 1921 1111
rect 1959 1108 1993 1111
rect 2031 1108 2065 1111
rect 2103 1108 2137 1111
rect 2175 1108 2209 1111
rect 2247 1108 2281 1111
rect 2387 1111 2419 1142
rect 2419 1111 2421 1142
rect 2459 1111 2487 1142
rect 2487 1111 2493 1142
rect 2531 1111 2555 1142
rect 2555 1111 2565 1142
rect 2603 1111 2623 1142
rect 2623 1111 2637 1142
rect 2675 1111 2691 1142
rect 2691 1111 2709 1142
rect 2747 1111 2759 1142
rect 2759 1111 2781 1142
rect 2819 1111 2827 1142
rect 2827 1111 2853 1142
rect 2891 1111 2895 1142
rect 2895 1111 2925 1142
rect 2963 1111 2997 1142
rect 3035 1111 3065 1142
rect 3065 1111 3069 1142
rect 3107 1111 3133 1142
rect 3133 1111 3141 1142
rect 3179 1111 3201 1142
rect 3201 1111 3213 1142
rect 2387 1108 2421 1111
rect 2459 1108 2493 1111
rect 2531 1108 2565 1111
rect 2603 1108 2637 1111
rect 2675 1108 2709 1111
rect 2747 1108 2781 1111
rect 2819 1108 2853 1111
rect 2891 1108 2925 1111
rect 2963 1108 2997 1111
rect 3035 1108 3069 1111
rect 3107 1108 3141 1111
rect 3179 1108 3213 1111
rect 3350 1111 3369 1142
rect 3369 1111 3384 1142
rect 3422 1111 3437 1142
rect 3437 1111 3456 1142
rect 3494 1111 3505 1142
rect 3505 1111 3528 1142
rect 3566 1111 3573 1142
rect 3573 1111 3600 1142
rect 3638 1111 3641 1142
rect 3641 1111 3672 1142
rect 3710 1111 3743 1142
rect 3743 1111 3744 1142
rect 3782 1111 3811 1142
rect 3811 1111 3816 1142
rect 3854 1111 3879 1142
rect 3879 1111 3888 1142
rect 3926 1111 3947 1142
rect 3947 1111 3960 1142
rect 3998 1111 4015 1142
rect 4015 1111 4032 1142
rect 4070 1111 4083 1142
rect 4083 1111 4104 1142
rect 4142 1111 4151 1142
rect 4151 1111 4176 1142
rect 4214 1111 4219 1142
rect 4219 1111 4248 1142
rect 4286 1111 4287 1142
rect 4287 1111 4320 1142
rect 4358 1111 4389 1142
rect 4389 1111 4392 1142
rect 4430 1111 4457 1142
rect 4457 1111 4464 1142
rect 4502 1111 4525 1142
rect 4525 1111 4536 1142
rect 4574 1111 4593 1142
rect 4593 1111 4608 1142
rect 4646 1111 4661 1142
rect 4661 1111 4680 1142
rect 4718 1111 4729 1142
rect 4729 1111 4752 1142
rect 4831 1111 4835 1142
rect 4835 1111 4865 1142
rect 4903 1111 4937 1142
rect 4975 1111 5005 1142
rect 5005 1111 5009 1142
rect 5047 1111 5073 1142
rect 5073 1111 5081 1142
rect 5119 1111 5141 1142
rect 5141 1111 5153 1142
rect 5191 1111 5209 1142
rect 5209 1111 5225 1142
rect 5263 1111 5277 1142
rect 5277 1111 5297 1142
rect 5335 1111 5345 1142
rect 5345 1111 5369 1142
rect 3350 1108 3384 1111
rect 3422 1108 3456 1111
rect 3494 1108 3528 1111
rect 3566 1108 3600 1111
rect 3638 1108 3672 1111
rect 3710 1108 3744 1111
rect 3782 1108 3816 1111
rect 3854 1108 3888 1111
rect 3926 1108 3960 1111
rect 3998 1108 4032 1111
rect 4070 1108 4104 1111
rect 4142 1108 4176 1111
rect 4214 1108 4248 1111
rect 4286 1108 4320 1111
rect 4358 1108 4392 1111
rect 4430 1108 4464 1111
rect 4502 1108 4536 1111
rect 4574 1108 4608 1111
rect 4646 1108 4680 1111
rect 4718 1108 4752 1111
rect 4831 1108 4865 1111
rect 4903 1108 4937 1111
rect 4975 1108 5009 1111
rect 5047 1108 5081 1111
rect 5119 1108 5153 1111
rect 5191 1108 5225 1111
rect 5263 1108 5297 1111
rect 5335 1108 5369 1111
rect 1175 1043 1209 1073
rect 1175 1039 1209 1043
rect 1289 1039 1304 1062
rect 1304 1039 1323 1062
rect 1361 1039 1373 1062
rect 1373 1039 1395 1062
rect 1433 1039 1442 1062
rect 1442 1039 1467 1062
rect 1505 1039 1511 1062
rect 1511 1039 1539 1062
rect 1577 1039 1580 1062
rect 1580 1039 1611 1062
rect 1649 1039 1683 1062
rect 1721 1039 1752 1062
rect 1752 1039 1755 1062
rect 1793 1039 1821 1062
rect 1821 1039 1827 1062
rect 1865 1039 1890 1062
rect 1890 1039 1899 1062
rect 1937 1039 1959 1062
rect 1959 1039 1971 1062
rect 2009 1039 2028 1062
rect 2028 1039 2043 1062
rect 2081 1039 2097 1062
rect 2097 1039 2115 1062
rect 2153 1039 2166 1062
rect 2166 1039 2187 1062
rect 2225 1039 2235 1062
rect 2235 1039 2259 1062
rect 2297 1039 2304 1062
rect 2304 1039 2331 1062
rect 2369 1039 2373 1062
rect 2373 1039 2403 1062
rect 2441 1039 2442 1062
rect 2442 1039 2475 1062
rect 2513 1039 2546 1062
rect 2546 1039 2547 1062
rect 2585 1039 2615 1062
rect 2615 1039 2619 1062
rect 2657 1039 2683 1062
rect 2683 1039 2691 1062
rect 2729 1039 2751 1062
rect 2751 1039 2763 1062
rect 2801 1039 2819 1062
rect 2819 1039 2835 1062
rect 1289 1028 1323 1039
rect 1361 1028 1395 1039
rect 1433 1028 1467 1039
rect 1505 1028 1539 1039
rect 1577 1028 1611 1039
rect 1649 1028 1683 1039
rect 1721 1028 1755 1039
rect 1793 1028 1827 1039
rect 1865 1028 1899 1039
rect 1937 1028 1971 1039
rect 2009 1028 2043 1039
rect 2081 1028 2115 1039
rect 2153 1028 2187 1039
rect 2225 1028 2259 1039
rect 2297 1028 2331 1039
rect 2369 1028 2403 1039
rect 2441 1028 2475 1039
rect 2513 1028 2547 1039
rect 2585 1028 2619 1039
rect 2657 1028 2691 1039
rect 2729 1028 2763 1039
rect 2801 1028 2835 1039
rect 3298 1039 3328 1062
rect 3328 1039 3332 1062
rect 3370 1039 3397 1062
rect 3397 1039 3404 1062
rect 3442 1039 3466 1062
rect 3466 1039 3476 1062
rect 3514 1039 3535 1062
rect 3535 1039 3548 1062
rect 3586 1039 3604 1062
rect 3604 1039 3620 1062
rect 3658 1039 3673 1062
rect 3673 1039 3692 1062
rect 3730 1039 3742 1062
rect 3742 1039 3764 1062
rect 3802 1039 3811 1062
rect 3811 1039 3836 1062
rect 3874 1039 3880 1062
rect 3880 1039 3908 1062
rect 3946 1039 3948 1062
rect 3948 1039 3980 1062
rect 4018 1039 4050 1062
rect 4050 1039 4052 1062
rect 4090 1039 4118 1062
rect 4118 1039 4124 1062
rect 4162 1039 4186 1062
rect 4186 1039 4196 1062
rect 4234 1039 4254 1062
rect 4254 1039 4268 1062
rect 4306 1039 4322 1062
rect 4322 1039 4340 1062
rect 4378 1039 4390 1062
rect 4390 1039 4412 1062
rect 4450 1039 4458 1062
rect 4458 1039 4484 1062
rect 4522 1039 4526 1062
rect 4526 1039 4556 1062
rect 3298 1028 3332 1039
rect 3370 1028 3404 1039
rect 3442 1028 3476 1039
rect 3514 1028 3548 1039
rect 3586 1028 3620 1039
rect 3658 1028 3692 1039
rect 3730 1028 3764 1039
rect 3802 1028 3836 1039
rect 3874 1028 3908 1039
rect 3946 1028 3980 1039
rect 4018 1028 4052 1039
rect 4090 1028 4124 1039
rect 4162 1028 4196 1039
rect 4234 1028 4268 1039
rect 4306 1028 4340 1039
rect 4378 1028 4412 1039
rect 4450 1028 4484 1039
rect 4522 1028 4556 1039
rect 1705 961 1739 988
rect 1777 961 1811 988
rect 1849 961 1883 988
rect 1921 961 1955 988
rect 1705 954 1717 961
rect 1717 954 1739 961
rect 1777 954 1785 961
rect 1785 954 1811 961
rect 1849 954 1853 961
rect 1853 954 1883 961
rect 1921 954 1955 961
rect 3563 927 3595 961
rect 3595 927 3597 961
rect 3635 927 3663 961
rect 3663 927 3669 961
rect 3707 927 3731 961
rect 3731 927 3741 961
rect 3779 927 3799 961
rect 3799 927 3813 961
rect 3851 927 3867 961
rect 3867 927 3885 961
rect 3923 927 3935 961
rect 3935 927 3957 961
rect 3995 927 4003 961
rect 4003 927 4029 961
rect 4067 927 4071 961
rect 4071 927 4101 961
rect 4139 927 4173 961
rect 4211 927 4241 961
rect 4241 927 4245 961
rect 4283 927 4309 961
rect 4309 927 4317 961
rect 5663 1039 5687 1062
rect 5687 1039 5697 1062
rect 5735 1039 5758 1062
rect 5758 1039 5769 1062
rect 5807 1039 5829 1062
rect 5829 1039 5841 1062
rect 5879 1039 5900 1062
rect 5900 1039 5913 1062
rect 5951 1039 5970 1062
rect 5970 1039 5985 1062
rect 5663 1028 5697 1039
rect 5735 1028 5769 1039
rect 5807 1028 5841 1039
rect 5879 1028 5913 1039
rect 5951 1028 5985 1039
rect 4978 927 4986 961
rect 4986 927 5012 961
rect 5050 927 5084 961
rect 5122 927 5156 961
rect 5194 927 5224 961
rect 5224 927 5228 961
rect 622 879 656 913
rect 694 879 728 913
rect 2048 879 2082 913
rect 2120 879 2154 913
rect 2192 879 2226 913
rect 2264 879 2298 913
rect 822 801 856 833
rect 822 799 856 801
rect 822 733 856 761
rect 822 727 856 733
rect 822 665 856 689
rect 822 655 856 665
rect 634 563 646 575
rect 646 563 668 575
rect 634 541 668 563
rect 634 461 668 495
rect 634 393 668 416
rect 634 382 646 393
rect 646 382 668 393
rect 822 597 856 611
rect 822 577 856 597
rect 822 495 856 528
rect 822 494 856 495
rect 822 427 856 446
rect 822 412 856 427
rect 634 325 668 337
rect 634 303 646 325
rect 646 303 668 325
rect 1174 801 1208 833
rect 1174 799 1208 801
rect 1174 733 1208 761
rect 1174 727 1208 733
rect 1174 665 1208 689
rect 1174 655 1208 665
rect 998 563 1032 575
rect 998 541 1032 563
rect 998 461 1032 495
rect 998 393 1032 416
rect 998 382 1032 393
rect 1174 597 1208 611
rect 1174 577 1208 597
rect 1174 495 1208 528
rect 1174 494 1208 495
rect 1174 427 1208 446
rect 1174 412 1208 427
rect 998 325 1032 337
rect 998 303 1032 325
rect 1526 801 1560 833
rect 1526 799 1560 801
rect 1526 733 1560 761
rect 1526 727 1560 733
rect 1526 665 1560 689
rect 1526 655 1560 665
rect 1350 563 1384 575
rect 1350 541 1384 563
rect 1350 461 1384 495
rect 1350 393 1384 416
rect 1350 382 1384 393
rect 1526 597 1560 611
rect 1526 577 1560 597
rect 1526 495 1560 528
rect 1526 494 1560 495
rect 1526 427 1560 446
rect 1526 412 1560 427
rect 1350 325 1384 337
rect 1350 303 1384 325
rect 1636 563 1670 596
rect 1636 562 1670 563
rect 1636 495 1670 504
rect 1636 470 1670 495
rect 1636 393 1670 413
rect 1636 379 1670 393
rect 1812 495 1846 516
rect 1812 482 1846 495
rect 1812 393 1846 426
rect 1812 392 1846 393
rect 1812 325 1846 337
rect 1812 303 1846 325
rect 1988 563 2022 596
rect 1988 562 2022 563
rect 1988 495 2022 509
rect 1988 475 2022 495
rect 1988 393 2022 423
rect 1988 389 2022 393
rect 1988 325 2022 337
rect 1988 303 2022 325
rect 2164 495 2198 516
rect 2164 482 2198 495
rect 2164 393 2198 426
rect 2164 392 2198 393
rect 2164 325 2198 337
rect 2164 303 2198 325
rect 2450 801 2484 833
rect 2450 799 2484 801
rect 2450 733 2484 761
rect 2450 727 2484 733
rect 2450 665 2484 689
rect 2450 655 2484 665
rect 2340 563 2374 596
rect 2340 562 2374 563
rect 2340 495 2374 509
rect 2340 475 2374 495
rect 2340 393 2374 423
rect 2340 389 2374 393
rect 2340 325 2374 337
rect 2340 303 2374 325
rect 2450 597 2484 611
rect 2450 577 2484 597
rect 2450 495 2484 526
rect 2450 492 2484 495
rect 2450 427 2484 441
rect 2450 407 2484 427
rect 2450 325 2484 357
rect 2450 323 2484 325
rect 2802 801 2836 833
rect 2802 799 2836 801
rect 2802 733 2836 761
rect 2802 727 2836 733
rect 2802 665 2836 689
rect 2802 655 2836 665
rect 2626 563 2660 596
rect 2626 562 2660 563
rect 2626 495 2660 509
rect 2626 475 2660 495
rect 2626 393 2660 423
rect 2626 389 2660 393
rect 2802 597 2836 611
rect 2802 577 2836 597
rect 2802 495 2836 528
rect 2802 494 2836 495
rect 2802 427 2836 445
rect 2802 411 2836 427
rect 2626 325 2660 337
rect 2626 303 2660 325
rect 3154 801 3188 833
rect 3154 799 3188 801
rect 3154 733 3188 761
rect 3154 727 3188 733
rect 3154 665 3188 689
rect 3154 655 3188 665
rect 2978 563 3012 596
rect 2978 562 3012 563
rect 2978 495 3012 509
rect 2978 475 3012 495
rect 2978 393 3012 423
rect 2978 389 3012 393
rect 3154 597 3188 611
rect 3154 577 3188 597
rect 3154 495 3188 528
rect 3154 494 3188 495
rect 3154 427 3188 445
rect 3154 411 3188 427
rect 2978 325 3012 337
rect 2978 303 3012 325
rect 3506 801 3540 833
rect 3506 799 3540 801
rect 3506 733 3540 761
rect 3506 727 3540 733
rect 3506 665 3540 689
rect 3506 655 3540 665
rect 3330 563 3364 596
rect 3330 562 3364 563
rect 3330 495 3364 509
rect 3330 475 3364 495
rect 3330 393 3364 423
rect 3330 389 3364 393
rect 3330 325 3364 337
rect 3330 303 3364 325
rect 3506 597 3540 611
rect 3506 577 3540 597
rect 3506 495 3540 521
rect 3506 487 3540 495
rect 3506 427 3540 431
rect 3506 397 3540 427
rect 3506 325 3540 341
rect 3506 307 3540 325
rect 3858 801 3892 833
rect 3858 799 3892 801
rect 3858 733 3892 761
rect 3858 727 3892 733
rect 3858 665 3892 689
rect 3858 655 3892 665
rect 3682 563 3716 596
rect 3682 562 3716 563
rect 3682 495 3716 509
rect 3682 475 3716 495
rect 3682 393 3716 423
rect 3682 389 3716 393
rect 3858 597 3892 611
rect 3858 577 3892 597
rect 3858 495 3892 528
rect 3858 494 3892 495
rect 3858 427 3892 445
rect 3858 411 3892 427
rect 3682 325 3716 337
rect 3682 303 3716 325
rect 4210 801 4244 833
rect 4210 799 4244 801
rect 4210 733 4244 761
rect 4210 727 4244 733
rect 4210 665 4244 689
rect 4210 655 4244 665
rect 4034 563 4068 596
rect 4034 562 4068 563
rect 4034 495 4068 509
rect 4034 475 4068 495
rect 4034 393 4068 423
rect 4034 389 4068 393
rect 4210 597 4244 611
rect 4210 577 4244 597
rect 4210 495 4244 528
rect 4210 494 4244 495
rect 4210 427 4244 445
rect 4210 411 4244 427
rect 4034 325 4068 337
rect 4034 303 4068 325
rect 4386 563 4420 596
rect 4386 562 4420 563
rect 4386 495 4420 509
rect 4386 475 4420 495
rect 4386 393 4420 423
rect 4386 389 4420 393
rect 4386 325 4420 337
rect 4386 303 4420 325
rect 4562 801 4596 833
rect 4562 799 4596 801
rect 4562 733 4596 761
rect 4562 727 4596 733
rect 4562 665 4596 689
rect 4562 655 4596 665
rect 4914 801 4948 833
rect 4914 799 4948 801
rect 4914 733 4948 761
rect 4914 727 4948 733
rect 4914 665 4948 689
rect 4914 655 4948 665
rect 4738 563 4772 596
rect 4738 562 4772 563
rect 4738 495 4772 509
rect 4738 475 4772 495
rect 4738 393 4772 423
rect 4738 389 4772 393
rect 4914 597 4948 611
rect 4914 577 4948 597
rect 4914 495 4948 528
rect 4914 494 4948 495
rect 4914 427 4948 445
rect 4914 411 4948 427
rect 4738 325 4772 337
rect 4738 303 4772 325
rect 5266 801 5300 833
rect 5266 799 5300 801
rect 5266 733 5300 761
rect 5266 727 5300 733
rect 5266 665 5300 689
rect 5266 655 5300 665
rect 5090 563 5124 596
rect 5090 562 5124 563
rect 5090 495 5124 509
rect 5090 475 5124 495
rect 5090 393 5124 423
rect 5090 389 5124 393
rect 5266 597 5300 611
rect 5266 577 5300 597
rect 5266 495 5300 528
rect 5266 494 5300 495
rect 5266 427 5300 445
rect 5266 411 5300 427
rect 5090 325 5124 337
rect 5090 303 5124 325
rect 5618 801 5652 833
rect 5618 799 5652 801
rect 5618 733 5652 761
rect 5618 727 5652 733
rect 5618 665 5652 689
rect 5618 655 5652 665
rect 5442 563 5476 596
rect 5442 562 5476 563
rect 5442 495 5476 509
rect 5442 475 5476 495
rect 5442 393 5476 423
rect 5442 389 5476 393
rect 5442 325 5476 337
rect 5442 303 5476 325
rect 5734 821 5768 833
rect 5734 799 5768 821
rect 5734 747 5768 761
rect 5734 727 5768 747
rect 5734 673 5768 689
rect 5734 655 5768 673
rect 5618 597 5652 611
rect 5618 577 5652 597
rect 5618 495 5652 521
rect 5618 487 5652 495
rect 5618 427 5652 431
rect 5618 397 5652 427
rect 5618 325 5652 341
rect 5618 307 5652 325
<< metal1 >>
rect 22 2223 6246 2235
rect 22 2189 88 2223
rect 122 2189 360 2223
rect 394 2189 802 2223
rect 836 2189 1114 2223
rect 1148 2189 1380 2223
rect 1414 2189 1692 2223
rect 1726 2189 2004 2223
rect 2038 2189 2316 2223
rect 2350 2189 2628 2223
rect 2662 2189 2940 2223
rect 2974 2189 3252 2223
rect 3286 2189 3604 2223
rect 3638 2189 3956 2223
rect 3990 2189 4308 2223
rect 4342 2189 4660 2223
rect 4694 2189 6134 2223
rect 6168 2189 6206 2223
rect 6240 2189 6246 2223
rect 22 2151 6246 2189
rect 22 2117 88 2151
rect 122 2117 360 2151
rect 394 2117 802 2151
rect 836 2117 1114 2151
rect 1148 2117 1380 2151
rect 1414 2117 1692 2151
rect 1726 2117 2004 2151
rect 2038 2117 2316 2151
rect 2350 2117 2628 2151
rect 2662 2117 2940 2151
rect 2974 2117 3252 2151
rect 3286 2117 3604 2151
rect 3638 2117 3956 2151
rect 3990 2117 4308 2151
rect 4342 2117 4660 2151
rect 4694 2117 6134 2151
rect 6168 2137 6246 2151
rect 6168 2117 6206 2137
rect 22 2103 6206 2117
rect 6240 2103 6246 2137
rect 22 2079 6246 2103
rect 22 2045 88 2079
rect 122 2045 360 2079
rect 394 2045 802 2079
rect 836 2045 1114 2079
rect 1148 2045 1380 2079
rect 1414 2045 1692 2079
rect 1726 2045 2004 2079
rect 2038 2045 2316 2079
rect 2350 2045 2628 2079
rect 2662 2045 2940 2079
rect 2974 2045 3252 2079
rect 3286 2045 3604 2079
rect 3638 2045 3956 2079
rect 3990 2045 4308 2079
rect 4342 2045 4660 2079
rect 4694 2045 6134 2079
rect 6168 2051 6246 2079
rect 6168 2045 6206 2051
rect 22 2033 6206 2045
rect -133 1998 388 2005
rect -133 1882 266 1998
rect 382 1882 388 1998
rect 1686 2001 1732 2033
rect -133 1875 388 1882
rect 1531 1974 1577 1986
rect 1531 1940 1537 1974
rect 1571 1940 1577 1974
rect 1531 1897 1577 1940
rect 1531 1863 1537 1897
rect 1571 1863 1577 1897
rect 1531 1820 1577 1863
rect 1531 1786 1537 1820
rect 1571 1786 1577 1820
rect 952 1741 998 1753
rect 952 1707 958 1741
rect 992 1707 998 1741
rect 952 1653 998 1707
rect 952 1619 958 1653
rect 992 1619 998 1653
rect 952 1572 998 1619
rect 1264 1741 1310 1753
rect 1264 1707 1270 1741
rect 1304 1707 1310 1741
rect 1264 1653 1310 1707
rect 1264 1619 1270 1653
rect 1304 1619 1310 1653
rect 1264 1572 1310 1619
rect 1531 1743 1577 1786
rect 1531 1709 1537 1743
rect 1571 1709 1577 1743
rect 1531 1666 1577 1709
rect 1531 1632 1537 1666
rect 1571 1632 1577 1666
rect 1686 1967 1692 2001
rect 1726 1967 1732 2001
rect 1998 2001 2044 2033
rect 1686 1925 1732 1967
rect 1686 1891 1692 1925
rect 1726 1891 1732 1925
rect 1686 1850 1732 1891
rect 1686 1816 1692 1850
rect 1726 1816 1732 1850
rect 1686 1775 1732 1816
rect 1686 1741 1692 1775
rect 1726 1741 1732 1775
rect 1686 1700 1732 1741
rect 1686 1666 1692 1700
rect 1726 1666 1732 1700
rect 1686 1634 1732 1666
rect 1842 1974 1888 1986
rect 1842 1940 1848 1974
rect 1882 1940 1888 1974
rect 1842 1897 1888 1940
rect 1842 1863 1848 1897
rect 1882 1863 1888 1897
rect 1842 1820 1888 1863
rect 1842 1786 1848 1820
rect 1882 1786 1888 1820
rect 1842 1743 1888 1786
rect 1842 1709 1848 1743
rect 1882 1709 1888 1743
rect 1842 1666 1888 1709
rect 1531 1595 1577 1632
rect 1842 1632 1848 1666
rect 1882 1632 1888 1666
rect 1998 1967 2004 2001
rect 2038 1967 2044 2001
rect 2310 2001 2356 2033
rect 1998 1925 2044 1967
rect 1998 1891 2004 1925
rect 2038 1891 2044 1925
rect 1998 1850 2044 1891
rect 1998 1816 2004 1850
rect 2038 1816 2044 1850
rect 1998 1775 2044 1816
rect 1998 1741 2004 1775
rect 2038 1741 2044 1775
rect 1998 1700 2044 1741
rect 1998 1666 2004 1700
rect 2038 1666 2044 1700
rect 1998 1634 2044 1666
rect 2154 1974 2200 1986
rect 2154 1940 2160 1974
rect 2194 1940 2200 1974
rect 2154 1897 2200 1940
rect 2154 1863 2160 1897
rect 2194 1863 2200 1897
rect 2154 1820 2200 1863
rect 2154 1786 2160 1820
rect 2194 1786 2200 1820
rect 2154 1743 2200 1786
rect 2154 1709 2160 1743
rect 2194 1709 2200 1743
rect 2154 1666 2200 1709
rect 1842 1595 1888 1632
rect 2154 1632 2160 1666
rect 2194 1632 2200 1666
rect 2310 1967 2316 2001
rect 2350 1967 2356 2001
rect 2310 1925 2356 1967
rect 2310 1891 2316 1925
rect 2350 1891 2356 1925
rect 2310 1850 2356 1891
rect 2310 1816 2316 1850
rect 2350 1816 2356 1850
rect 2310 1775 2356 1816
rect 2310 1741 2316 1775
rect 2350 1741 2356 1775
rect 2310 1700 2356 1741
rect 2310 1666 2316 1700
rect 2350 1666 2356 1700
rect 2622 2001 2668 2033
rect 2622 1967 2628 2001
rect 2662 1967 2668 2001
rect 2622 1923 2668 1967
rect 2934 2001 2980 2033
rect 2934 1967 2940 2001
rect 2974 1967 2980 2001
rect 2622 1889 2628 1923
rect 2662 1889 2668 1923
rect 2622 1845 2668 1889
rect 2622 1811 2628 1845
rect 2662 1811 2668 1845
rect 2622 1767 2668 1811
rect 2622 1733 2628 1767
rect 2662 1733 2668 1767
rect 2310 1634 2356 1666
rect 2539 1665 2591 1694
rect 2154 1595 2200 1632
rect 2539 1601 2591 1613
rect 1486 1589 2539 1595
rect 952 1566 1315 1572
rect 952 1532 958 1566
rect 992 1532 1270 1566
rect 1304 1532 1315 1566
rect 1486 1555 1537 1589
rect 1571 1555 1848 1589
rect 1882 1555 2160 1589
rect 2194 1555 2539 1589
rect 1486 1549 2539 1555
rect 1486 1543 2591 1549
rect 2622 1690 2668 1733
rect 2622 1656 2628 1690
rect 2662 1656 2668 1690
rect 2622 1613 2668 1656
rect 2622 1579 2628 1613
rect 2662 1579 2668 1613
rect 2622 1547 2668 1579
rect 2778 1939 2824 1951
rect 2778 1905 2784 1939
rect 2818 1905 2824 1939
rect 2778 1862 2824 1905
rect 2778 1828 2784 1862
rect 2818 1828 2824 1862
rect 2778 1785 2824 1828
rect 2778 1751 2784 1785
rect 2818 1751 2824 1785
rect 2778 1708 2824 1751
rect 2778 1674 2784 1708
rect 2818 1674 2824 1708
rect 2778 1632 2824 1674
rect 2778 1598 2784 1632
rect 2818 1598 2824 1632
rect 2934 1921 2980 1967
rect 3246 2001 3292 2033
rect 3246 1967 3252 2001
rect 3286 1967 3292 2001
rect 2934 1887 2940 1921
rect 2974 1887 2980 1921
rect 2934 1842 2980 1887
rect 2934 1808 2940 1842
rect 2974 1808 2980 1842
rect 2934 1763 2980 1808
rect 2934 1729 2940 1763
rect 2974 1729 2980 1763
rect 2934 1684 2980 1729
rect 2934 1650 2940 1684
rect 2974 1650 2980 1684
rect 2934 1618 2980 1650
rect 3091 1939 3137 1951
rect 3091 1905 3097 1939
rect 3131 1905 3137 1939
rect 3091 1862 3137 1905
rect 3091 1828 3097 1862
rect 3131 1828 3137 1862
rect 3091 1785 3137 1828
rect 3091 1751 3097 1785
rect 3131 1751 3137 1785
rect 3091 1708 3137 1751
rect 3091 1674 3097 1708
rect 3131 1674 3137 1708
rect 3091 1632 3137 1674
rect 2778 1556 2824 1598
rect 3091 1598 3097 1632
rect 3131 1598 3137 1632
rect 3246 1921 3292 1967
rect 3598 2001 3644 2033
rect 3598 1967 3604 2001
rect 3638 1967 3644 2001
rect 3246 1887 3252 1921
rect 3286 1887 3292 1921
rect 3246 1842 3292 1887
rect 3246 1808 3252 1842
rect 3286 1808 3292 1842
rect 3246 1763 3292 1808
rect 3246 1729 3252 1763
rect 3286 1729 3292 1763
rect 3246 1684 3292 1729
rect 3246 1650 3252 1684
rect 3286 1650 3292 1684
rect 3246 1618 3292 1650
rect 3422 1950 3468 1962
rect 3422 1916 3428 1950
rect 3462 1916 3468 1950
rect 3422 1873 3468 1916
rect 3422 1839 3428 1873
rect 3462 1839 3468 1873
rect 3422 1796 3468 1839
rect 3422 1762 3428 1796
rect 3462 1762 3468 1796
rect 3422 1719 3468 1762
rect 3422 1685 3428 1719
rect 3462 1685 3468 1719
rect 3422 1643 3468 1685
rect 3091 1559 3137 1598
rect 2991 1556 2997 1559
tri 2740 1547 2749 1556 se
rect 2749 1547 2784 1556
tri 2736 1543 2740 1547 se
rect 2740 1543 2784 1547
rect 952 1520 1315 1532
tri 2715 1522 2736 1543 se
rect 2736 1522 2784 1543
rect 2818 1522 2997 1556
tri 2714 1521 2715 1522 se
rect 2715 1521 2997 1522
tri 2713 1520 2714 1521 se
rect 2714 1520 2997 1521
tri 2687 1494 2713 1520 se
rect 2713 1510 2997 1520
rect 2713 1494 2770 1510
tri 2770 1494 2786 1510 nw
rect 2991 1507 2997 1510
rect 3049 1507 3061 1559
rect 3113 1556 3137 1559
rect 3422 1609 3428 1643
rect 3462 1609 3468 1643
rect 3598 1921 3644 1967
rect 3950 2001 3996 2033
rect 3950 1967 3956 2001
rect 3990 1967 3996 2001
rect 3598 1887 3604 1921
rect 3638 1887 3644 1921
rect 3598 1842 3644 1887
rect 3598 1808 3604 1842
rect 3638 1808 3644 1842
rect 3598 1763 3644 1808
rect 3598 1729 3604 1763
rect 3638 1729 3644 1763
rect 3598 1684 3644 1729
rect 3598 1650 3604 1684
rect 3638 1650 3644 1684
rect 3598 1618 3644 1650
rect 3774 1950 3820 1962
rect 3774 1916 3780 1950
rect 3814 1916 3820 1950
rect 3774 1873 3820 1916
rect 3774 1839 3780 1873
rect 3814 1839 3820 1873
rect 3774 1796 3820 1839
rect 3774 1762 3780 1796
rect 3814 1762 3820 1796
rect 3774 1719 3820 1762
rect 3774 1685 3780 1719
rect 3814 1685 3820 1719
rect 3774 1643 3820 1685
rect 3422 1567 3468 1609
rect 3774 1609 3780 1643
rect 3814 1609 3820 1643
rect 3950 1921 3996 1967
rect 4302 2001 4348 2033
rect 4302 1967 4308 2001
rect 4342 1967 4348 2001
rect 3950 1887 3956 1921
rect 3990 1887 3996 1921
rect 3950 1842 3996 1887
rect 3950 1808 3956 1842
rect 3990 1808 3996 1842
rect 3950 1763 3996 1808
rect 3950 1729 3956 1763
rect 3990 1729 3996 1763
rect 3950 1684 3996 1729
rect 3950 1650 3956 1684
rect 3990 1650 3996 1684
rect 3950 1618 3996 1650
rect 4126 1950 4172 1962
rect 4126 1916 4132 1950
rect 4166 1916 4172 1950
rect 4126 1873 4172 1916
rect 4126 1839 4132 1873
rect 4166 1839 4172 1873
rect 4126 1796 4172 1839
rect 4126 1762 4132 1796
rect 4166 1762 4172 1796
rect 4126 1719 4172 1762
rect 4126 1685 4132 1719
rect 4166 1685 4172 1719
rect 4126 1643 4172 1685
rect 3774 1567 3820 1609
rect 4126 1609 4132 1643
rect 4166 1609 4172 1643
rect 4302 1921 4348 1967
rect 4654 2001 4700 2033
rect 4654 1967 4660 2001
rect 4694 1967 4700 2001
rect 6200 2017 6206 2033
rect 6240 2017 6246 2051
rect 4302 1887 4308 1921
rect 4342 1887 4348 1921
rect 4302 1842 4348 1887
rect 4302 1808 4308 1842
rect 4342 1808 4348 1842
rect 4302 1763 4348 1808
rect 4302 1729 4308 1763
rect 4342 1729 4348 1763
rect 4302 1684 4348 1729
rect 4302 1650 4308 1684
rect 4342 1650 4348 1684
rect 4302 1618 4348 1650
rect 4478 1950 4524 1962
rect 4478 1916 4484 1950
rect 4518 1916 4524 1950
rect 4478 1873 4524 1916
rect 4478 1839 4484 1873
rect 4518 1839 4524 1873
rect 4478 1796 4524 1839
rect 4478 1762 4484 1796
rect 4518 1762 4524 1796
rect 4478 1719 4524 1762
rect 4478 1685 4484 1719
rect 4518 1685 4524 1719
rect 4478 1643 4524 1685
rect 4126 1567 4172 1609
rect 4478 1609 4484 1643
rect 4518 1609 4524 1643
rect 4654 1921 4700 1967
rect 4654 1887 4660 1921
rect 4694 1887 4700 1921
rect 4654 1842 4700 1887
rect 4654 1808 4660 1842
rect 4694 1808 4700 1842
rect 4654 1763 4700 1808
rect 4654 1729 4660 1763
rect 4694 1729 4700 1763
rect 4654 1684 4700 1729
rect 4654 1650 4660 1684
rect 4694 1650 4700 1684
rect 4654 1618 4700 1650
rect 4764 1973 6058 1985
rect 4764 1939 4770 1973
rect 4804 1939 5082 1973
rect 5116 1939 5394 1973
rect 5428 1939 5706 1973
rect 5740 1939 6018 1973
rect 6052 1939 6058 1973
rect 4764 1891 4810 1939
rect 4764 1857 4770 1891
rect 4804 1857 4810 1891
rect 5076 1891 5122 1939
rect 4764 1809 4810 1857
rect 4764 1775 4770 1809
rect 4804 1775 4810 1809
rect 4764 1728 4810 1775
rect 4764 1694 4770 1728
rect 4804 1694 4810 1728
rect 4764 1647 4810 1694
rect 4478 1567 4524 1609
rect 4764 1613 4770 1647
rect 4804 1613 4810 1647
rect 4764 1601 4810 1613
rect 4920 1869 4966 1881
rect 4920 1835 4926 1869
rect 4960 1835 4966 1869
rect 4920 1793 4966 1835
rect 4920 1759 4926 1793
rect 4960 1759 4966 1793
rect 4920 1717 4966 1759
rect 4920 1683 4926 1717
rect 4960 1683 4966 1717
rect 4920 1642 4966 1683
rect 4920 1608 4926 1642
rect 4960 1608 4966 1642
rect 4920 1567 4966 1608
rect 5076 1857 5082 1891
rect 5116 1857 5122 1891
rect 5388 1897 5434 1939
rect 5076 1809 5122 1857
rect 5076 1775 5082 1809
rect 5116 1775 5122 1809
rect 5076 1728 5122 1775
rect 5076 1694 5082 1728
rect 5116 1694 5122 1728
rect 5076 1647 5122 1694
rect 5076 1613 5082 1647
rect 5116 1613 5122 1647
rect 5076 1601 5122 1613
rect 5233 1869 5279 1881
rect 5233 1835 5239 1869
rect 5273 1835 5279 1869
rect 5233 1783 5279 1835
rect 5233 1749 5239 1783
rect 5273 1749 5279 1783
rect 5233 1698 5279 1749
rect 5233 1664 5239 1698
rect 5273 1664 5279 1698
rect 5233 1613 5279 1664
rect 5233 1579 5239 1613
rect 5273 1579 5279 1613
rect 5233 1567 5279 1579
rect 3131 1522 3142 1556
rect 3113 1510 3142 1522
rect 3422 1533 3428 1567
rect 3462 1533 3780 1567
rect 3814 1533 4132 1567
rect 4166 1533 4484 1567
rect 4518 1533 4926 1567
rect 4960 1533 5279 1567
rect 3422 1528 5279 1533
rect 3422 1521 5239 1528
rect 3113 1507 3119 1510
rect 5233 1494 5239 1521
rect 5273 1494 5279 1528
tri 2677 1484 2687 1494 se
rect 2687 1484 2760 1494
tri 2760 1484 2770 1494 nw
rect 1163 1432 1169 1484
rect 1221 1432 1233 1484
rect 1285 1478 2335 1484
tri 2335 1478 2341 1484 sw
tri 2672 1479 2677 1484 se
rect 2677 1479 2754 1484
rect 2413 1478 2565 1479
tri 2671 1478 2672 1479 se
rect 2672 1478 2754 1479
tri 2754 1478 2760 1484 nw
rect 1285 1473 2735 1478
rect 1285 1439 2425 1473
rect 2459 1439 2519 1473
rect 2553 1459 2735 1473
tri 2735 1459 2754 1478 nw
rect 2553 1447 2723 1459
tri 2723 1447 2735 1459 nw
rect 2553 1443 2719 1447
tri 2719 1443 2723 1447 nw
rect 2553 1439 2708 1443
rect 1285 1432 2708 1439
tri 2708 1432 2719 1443 nw
rect 2817 1425 2823 1477
rect 2875 1425 2887 1477
rect 2939 1425 4572 1477
rect 4624 1425 4636 1477
rect 4688 1459 5092 1477
tri 5092 1459 5110 1477 sw
rect 4688 1447 5110 1459
tri 5110 1447 5122 1459 sw
rect 4688 1443 5122 1447
tri 5122 1443 5126 1447 sw
rect 5233 1443 5279 1494
rect 4688 1432 5126 1443
tri 5126 1432 5137 1443 sw
rect 4688 1426 5137 1432
tri 5137 1426 5143 1432 sw
rect 4688 1425 5143 1426
tri 5061 1409 5077 1425 ne
rect 5077 1409 5143 1425
tri 5143 1409 5160 1426 sw
rect 5233 1409 5239 1443
rect 5273 1409 5279 1443
tri 5077 1381 5105 1409 ne
rect 5105 1397 5160 1409
tri 5160 1397 5172 1409 sw
rect 5233 1397 5279 1409
rect 5388 1863 5394 1897
rect 5428 1863 5434 1897
rect 5388 1821 5434 1863
rect 5388 1787 5394 1821
rect 5428 1787 5434 1821
rect 5388 1745 5434 1787
rect 5388 1711 5394 1745
rect 5428 1711 5434 1745
rect 5388 1669 5434 1711
rect 5388 1635 5394 1669
rect 5428 1635 5434 1669
rect 5388 1593 5434 1635
rect 5388 1559 5394 1593
rect 5428 1559 5434 1593
rect 5388 1518 5434 1559
rect 5388 1484 5394 1518
rect 5428 1484 5434 1518
rect 5388 1443 5434 1484
rect 5388 1409 5394 1443
rect 5428 1409 5434 1443
rect 5388 1397 5434 1409
rect 5544 1887 5590 1899
rect 5544 1853 5550 1887
rect 5584 1853 5590 1887
rect 5544 1808 5590 1853
rect 5544 1774 5550 1808
rect 5584 1774 5590 1808
rect 5544 1729 5590 1774
rect 5544 1695 5550 1729
rect 5584 1695 5590 1729
rect 5544 1650 5590 1695
rect 5544 1616 5550 1650
rect 5584 1616 5590 1650
rect 5544 1571 5590 1616
rect 5544 1537 5550 1571
rect 5584 1537 5590 1571
rect 5544 1493 5590 1537
rect 5544 1459 5550 1493
rect 5584 1459 5590 1493
rect 5544 1415 5590 1459
rect 5105 1381 5172 1397
tri 5172 1381 5188 1397 sw
rect 5544 1381 5550 1415
rect 5584 1381 5590 1415
rect 5700 1897 5746 1939
rect 5700 1863 5706 1897
rect 5740 1863 5746 1897
rect 5700 1821 5746 1863
rect 5700 1787 5706 1821
rect 5740 1787 5746 1821
rect 5700 1745 5746 1787
rect 5700 1711 5706 1745
rect 5740 1711 5746 1745
rect 5700 1669 5746 1711
rect 5700 1635 5706 1669
rect 5740 1635 5746 1669
rect 5700 1593 5746 1635
rect 5700 1559 5706 1593
rect 5740 1559 5746 1593
rect 5700 1518 5746 1559
rect 5700 1484 5706 1518
rect 5740 1484 5746 1518
rect 5700 1443 5746 1484
rect 5700 1409 5706 1443
rect 5740 1409 5746 1443
rect 5700 1397 5746 1409
rect 5856 1887 5902 1899
rect 5856 1853 5862 1887
rect 5896 1853 5902 1887
rect 5856 1808 5902 1853
rect 5856 1774 5862 1808
rect 5896 1774 5902 1808
rect 5856 1729 5902 1774
rect 5856 1695 5862 1729
rect 5896 1695 5902 1729
rect 5856 1650 5902 1695
rect 5856 1616 5862 1650
rect 5896 1616 5902 1650
rect 5856 1572 5902 1616
rect 5856 1538 5862 1572
rect 5896 1538 5902 1572
rect 5856 1494 5902 1538
rect 5856 1460 5862 1494
rect 5896 1460 5902 1494
rect 5856 1416 5902 1460
tri 5105 1365 5121 1381 ne
rect 5121 1365 5188 1381
tri 5188 1365 5204 1381 sw
tri 5121 1343 5143 1365 ne
rect 5143 1343 5204 1365
tri 5204 1343 5226 1365 sw
rect 5544 1343 5590 1381
rect 5856 1382 5862 1416
rect 5896 1382 5902 1416
rect 5856 1343 5902 1382
tri 5143 1340 5146 1343 ne
rect 5146 1340 5902 1343
tri 5146 1338 5148 1340 ne
rect 5148 1338 5902 1340
tri 5148 1337 5149 1338 ne
rect 5149 1337 5862 1338
tri 5149 1303 5183 1337 ne
rect 5183 1303 5550 1337
rect 5584 1304 5862 1337
rect 5896 1304 5902 1338
rect 5584 1303 5902 1304
tri 5183 1294 5192 1303 ne
rect 5192 1294 5902 1303
rect 6012 1893 6058 1939
rect 6012 1859 6018 1893
rect 6052 1859 6058 1893
rect 6012 1814 6058 1859
rect 6012 1780 6018 1814
rect 6052 1780 6058 1814
rect 6200 1965 6246 2017
rect 6200 1931 6206 1965
rect 6240 1931 6246 1965
rect 6200 1879 6246 1931
rect 6200 1845 6206 1879
rect 6240 1845 6246 1879
rect 6200 1813 6246 1845
rect 6012 1735 6058 1780
rect 6012 1701 6018 1735
rect 6052 1701 6058 1735
rect 6012 1656 6058 1701
rect 6012 1622 6018 1656
rect 6052 1622 6058 1656
rect 6012 1577 6058 1622
rect 6012 1543 6018 1577
rect 6052 1543 6058 1577
rect 6012 1498 6058 1543
rect 6012 1464 6018 1498
rect 6052 1464 6058 1498
rect 6012 1419 6058 1464
rect 6012 1385 6018 1419
rect 6052 1385 6058 1419
rect 6012 1340 6058 1385
rect 6128 1767 6246 1813
rect 6128 1726 6174 1767
rect 6128 1692 6134 1726
rect 6168 1692 6174 1726
rect 6128 1645 6174 1692
rect 6128 1611 6134 1645
rect 6168 1611 6174 1645
rect 6128 1563 6174 1611
rect 6128 1529 6134 1563
rect 6168 1529 6174 1563
rect 6128 1481 6174 1529
rect 6128 1447 6134 1481
rect 6168 1447 6174 1481
rect 6128 1399 6174 1447
rect 6128 1365 6134 1399
rect 6168 1365 6174 1399
rect 6128 1363 6174 1365
rect 6012 1306 6018 1340
rect 6052 1306 6058 1340
rect 6012 1294 6058 1306
rect 6122 1357 6174 1363
tri 5192 1291 5195 1294 ne
rect 5195 1292 5902 1294
rect 5195 1291 5901 1292
rect 6122 1283 6134 1305
rect 6168 1283 6174 1305
rect 6122 1247 6174 1283
rect 452 1228 4764 1240
rect 452 1194 464 1228
rect 498 1194 536 1228
rect 570 1194 4764 1228
rect 452 1188 4764 1194
rect 6122 1189 6174 1195
tri 3313 1163 3338 1188 ne
rect 184 1154 930 1160
rect 184 1120 196 1154
rect 230 1120 268 1154
rect 302 1120 340 1154
rect 374 1120 412 1154
rect 446 1145 930 1154
rect 446 1120 890 1145
rect 184 1114 890 1120
tri 859 1111 862 1114 ne
rect 862 1111 890 1114
rect 924 1111 930 1145
tri 862 1108 865 1111 ne
rect 865 1108 930 1111
tri 865 1096 877 1108 ne
rect 877 1096 930 1108
tri 877 1089 884 1096 ne
rect -47 1073 62 1086
tri 62 1073 75 1086 sw
rect 884 1073 930 1096
rect -47 1068 75 1073
tri 75 1068 80 1073 sw
rect -47 1039 80 1068
tri 80 1039 109 1068 sw
rect 884 1039 890 1073
rect 924 1039 930 1073
rect -47 1028 109 1039
tri 109 1028 120 1039 sw
rect -47 1027 120 1028
tri 120 1027 121 1028 sw
rect 884 1027 930 1039
rect 1030 1145 1076 1157
rect 1030 1111 1036 1145
rect 1070 1111 1076 1145
rect 1030 1073 1076 1111
rect 1030 1039 1036 1073
rect 1070 1039 1076 1073
rect -47 988 121 1027
tri 121 988 160 1027 sw
rect -47 954 160 988
tri 160 954 194 988 sw
rect -47 944 194 954
tri 194 944 204 954 sw
rect -47 927 204 944
tri 204 927 221 944 sw
tri 1013 927 1030 944 se
rect 1030 927 1076 1039
rect 1163 1151 1215 1157
rect 1163 1087 1215 1099
rect 1443 1142 2124 1148
rect 2176 1142 2188 1148
rect 2240 1142 2293 1148
rect 1443 1108 1455 1142
rect 1489 1108 1527 1142
rect 1561 1108 1599 1142
rect 1633 1108 1671 1142
rect 1705 1108 1743 1142
rect 1777 1108 1815 1142
rect 1849 1108 1887 1142
rect 1921 1108 1959 1142
rect 1993 1108 2031 1142
rect 2065 1108 2103 1142
rect 2240 1108 2247 1142
rect 2281 1108 2293 1142
rect 1443 1096 2124 1108
rect 2176 1096 2188 1108
rect 2240 1096 2293 1108
rect 2375 1142 2823 1148
rect 2375 1108 2387 1142
rect 2421 1108 2459 1142
rect 2493 1108 2531 1142
rect 2565 1108 2603 1142
rect 2637 1108 2675 1142
rect 2709 1108 2747 1142
rect 2781 1108 2819 1142
rect 2375 1096 2823 1108
rect 2875 1096 2887 1148
rect 2939 1142 3225 1148
rect 2939 1108 2963 1142
rect 2997 1108 3035 1142
rect 3069 1108 3107 1142
rect 3141 1108 3179 1142
rect 3213 1108 3225 1142
rect 2939 1096 3225 1108
rect 3338 1142 4764 1188
tri 6194 1148 6202 1156 se
rect 6202 1148 6328 1156
rect 3338 1108 3350 1142
rect 3384 1108 3422 1142
rect 3456 1108 3494 1142
rect 3528 1108 3566 1142
rect 3600 1108 3638 1142
rect 3672 1108 3710 1142
rect 3744 1108 3782 1142
rect 3816 1108 3854 1142
rect 3888 1108 3926 1142
rect 3960 1108 3998 1142
rect 4032 1108 4070 1142
rect 4104 1108 4142 1142
rect 4176 1108 4214 1142
rect 4248 1108 4286 1142
rect 4320 1108 4358 1142
rect 4392 1108 4430 1142
rect 4464 1108 4502 1142
rect 4536 1108 4574 1142
rect 4608 1108 4646 1142
rect 4680 1108 4718 1142
rect 4752 1108 4764 1142
rect 3338 1096 4764 1108
rect 4819 1142 4982 1148
rect 4819 1108 4831 1142
rect 4865 1108 4903 1142
rect 4937 1108 4975 1142
rect 4819 1096 4982 1108
rect 5034 1096 5046 1148
rect 5098 1142 5381 1148
rect 5098 1108 5119 1142
rect 5153 1108 5191 1142
rect 5225 1108 5263 1142
rect 5297 1108 5335 1142
rect 5369 1108 5381 1142
rect 5098 1096 5381 1108
tri 6142 1096 6194 1148 se
rect 6194 1096 6328 1148
tri 6135 1089 6142 1096 se
rect 6142 1089 6328 1096
tri 6114 1068 6135 1089 se
rect 6135 1068 6328 1089
rect 1163 1023 1215 1035
rect 1277 1062 5770 1068
rect 5822 1062 5880 1068
rect 5932 1062 5997 1068
rect 1277 1028 1289 1062
rect 1323 1028 1361 1062
rect 1395 1028 1433 1062
rect 1467 1028 1505 1062
rect 1539 1028 1577 1062
rect 1611 1028 1649 1062
rect 1683 1028 1721 1062
rect 1755 1028 1793 1062
rect 1827 1028 1865 1062
rect 1899 1028 1937 1062
rect 1971 1028 2009 1062
rect 2043 1028 2081 1062
rect 2115 1028 2153 1062
rect 2187 1028 2225 1062
rect 2259 1028 2297 1062
rect 2331 1028 2369 1062
rect 2403 1028 2441 1062
rect 2475 1028 2513 1062
rect 2547 1028 2585 1062
rect 2619 1028 2657 1062
rect 2691 1028 2729 1062
rect 2763 1028 2801 1062
rect 2835 1028 3298 1062
rect 3332 1028 3370 1062
rect 3404 1028 3442 1062
rect 3476 1028 3514 1062
rect 3548 1028 3586 1062
rect 3620 1028 3658 1062
rect 3692 1028 3730 1062
rect 3764 1028 3802 1062
rect 3836 1028 3874 1062
rect 3908 1028 3946 1062
rect 3980 1028 4018 1062
rect 4052 1028 4090 1062
rect 4124 1028 4162 1062
rect 4196 1028 4234 1062
rect 4268 1028 4306 1062
rect 4340 1028 4378 1062
rect 4412 1028 4450 1062
rect 4484 1028 4522 1062
rect 4556 1028 5663 1062
rect 5697 1028 5735 1062
rect 5769 1028 5770 1062
rect 5841 1028 5879 1062
rect 5932 1028 5951 1062
rect 5985 1028 5997 1062
rect 1277 1022 5770 1028
tri 1215 994 1240 1019 sw
rect 5764 1016 5770 1022
rect 5822 1016 5880 1028
rect 5932 1022 5997 1028
tri 6068 1022 6114 1068 se
rect 6114 1022 6328 1068
rect 5932 1016 5938 1022
tri 6065 1019 6068 1022 se
rect 6068 1019 6328 1022
tri 6062 1016 6065 1019 se
rect 6065 1016 6328 1019
tri 6040 994 6062 1016 se
rect 6062 994 6328 1016
rect 1215 988 1967 994
rect 1215 971 1705 988
rect 1163 954 1705 971
rect 1739 954 1777 988
rect 1811 954 1849 988
rect 1883 954 1921 988
rect 1955 954 1967 988
tri 6013 967 6040 994 se
rect 6040 967 6328 994
rect 1163 948 1967 954
tri 1076 927 1093 944 sw
rect -47 919 221 927
tri 221 919 229 927 sw
tri 1005 919 1013 927 se
rect 1013 919 1093 927
tri 1093 919 1101 927 sw
rect -47 913 229 919
tri 229 913 235 919 sw
rect 610 913 2310 919
rect 2340 915 2346 967
rect 2398 915 2410 967
rect 2462 961 4343 967
rect 2462 927 3563 961
rect 3597 927 3635 961
rect 3669 927 3707 961
rect 3741 927 3779 961
rect 3813 927 3851 961
rect 3885 927 3923 961
rect 3957 927 3995 961
rect 4029 927 4067 961
rect 4101 927 4139 961
rect 4173 927 4211 961
rect 4245 927 4283 961
rect 4317 927 4343 961
rect 2462 915 4343 927
rect 4387 915 4393 967
rect 4445 915 4457 967
rect 4509 961 4982 967
rect 4509 927 4978 961
rect 4509 915 4982 927
rect 5034 915 5046 967
rect 5098 961 5240 967
rect 5098 927 5122 961
rect 5156 927 5194 961
rect 5228 927 5240 961
rect 5098 915 5240 927
tri 5961 915 6013 967 se
rect 6013 915 6328 967
rect -47 884 235 913
tri -47 879 -42 884 ne
rect -42 879 235 884
tri 235 879 269 913 sw
rect 610 879 622 913
rect 656 879 694 913
rect 728 879 2048 913
rect 2082 879 2120 913
rect 2154 879 2192 913
rect 2226 879 2264 913
rect 2298 879 2310 913
tri -42 845 -8 879 ne
rect -8 873 269 879
tri 269 873 275 879 sw
rect 610 873 2310 879
tri 5919 873 5961 915 se
rect 5961 873 6328 915
rect -8 845 275 873
tri 275 845 303 873 sw
tri 5891 845 5919 873 se
rect 5919 845 6328 873
tri -8 833 4 845 ne
rect 4 833 6328 845
tri 4 799 38 833 ne
rect 38 799 266 833
rect 394 799 822 833
rect 856 799 1174 833
rect 1208 799 1526 833
rect 1560 799 2450 833
rect 2484 799 2802 833
rect 2836 799 3154 833
rect 3188 799 3506 833
rect 3540 799 3858 833
rect 3892 799 4210 833
rect 4244 799 4562 833
rect 4596 799 4914 833
rect 4948 799 5266 833
rect 5300 799 5618 833
rect 5652 799 5734 833
rect 5768 799 6328 833
tri 38 775 62 799 ne
rect 62 775 266 799
tri 62 761 76 775 ne
rect 76 761 266 775
rect 382 761 6328 799
tri 76 740 97 761 ne
rect 97 740 266 761
rect -133 734 19 740
rect -133 484 -99 734
rect 7 611 19 734
tri 97 727 110 740 ne
rect 110 727 266 740
rect 394 727 822 761
rect 856 727 1174 761
rect 1208 727 1526 761
rect 1560 727 2450 761
rect 2484 727 2802 761
rect 2836 727 3154 761
rect 3188 727 3506 761
rect 3540 727 3858 761
rect 3892 727 4210 761
rect 4244 727 4562 761
rect 4596 727 4914 761
rect 4948 727 5266 761
rect 5300 727 5618 761
rect 5652 727 5734 761
rect 5768 727 6328 761
tri 110 689 148 727 ne
rect 148 689 266 727
rect 382 689 6328 727
tri 148 655 182 689 ne
rect 182 655 266 689
rect 394 655 822 689
rect 856 655 1174 689
rect 1208 655 1526 689
rect 1560 655 2450 689
rect 2484 655 2802 689
rect 2836 655 3154 689
rect 3188 655 3506 689
rect 3540 655 3858 689
rect 3892 655 4210 689
rect 4244 655 4562 689
rect 4596 655 4914 689
rect 4948 655 5266 689
rect 5300 655 5618 689
rect 5652 655 5734 689
rect 5768 655 6328 689
tri 182 643 194 655 ne
rect 194 653 266 655
rect 382 653 6328 655
rect 194 643 6328 653
tri 19 611 27 619 sw
rect 816 611 862 643
rect 7 594 27 611
tri 27 594 44 611 sw
rect 7 484 266 594
rect -133 478 266 484
rect 382 478 388 594
rect 628 575 674 587
rect 628 541 634 575
rect 668 541 674 575
rect 628 495 674 541
rect 628 461 634 495
rect 668 461 674 495
rect 628 416 674 461
rect 628 382 634 416
rect 668 382 674 416
rect 628 337 674 382
rect 816 577 822 611
rect 856 577 862 611
rect 1168 611 1214 643
rect 816 528 862 577
rect 816 494 822 528
rect 856 494 862 528
rect 816 446 862 494
rect 816 412 822 446
rect 856 412 862 446
rect 816 380 862 412
rect 992 575 1038 587
rect 992 541 998 575
rect 1032 541 1038 575
rect 992 495 1038 541
rect 992 461 998 495
rect 1032 461 1038 495
rect 992 416 1038 461
rect 992 382 998 416
rect 1032 382 1038 416
rect 628 303 634 337
rect 668 303 674 337
rect 628 291 674 303
rect 992 337 1038 382
rect 1168 577 1174 611
rect 1208 577 1214 611
rect 1520 611 1566 643
rect 1168 528 1214 577
rect 1168 494 1174 528
rect 1208 494 1214 528
rect 1168 446 1214 494
rect 1168 412 1174 446
rect 1208 412 1214 446
rect 1168 380 1214 412
rect 1344 575 1390 587
rect 1344 541 1350 575
rect 1384 541 1390 575
rect 1344 495 1390 541
rect 1344 461 1350 495
rect 1384 461 1390 495
rect 1344 416 1390 461
rect 1344 382 1350 416
rect 1384 382 1390 416
rect 1344 337 1390 382
rect 1520 577 1526 611
rect 1560 577 1566 611
rect 2444 611 2490 643
rect 1520 528 1566 577
rect 1520 494 1526 528
rect 1560 494 1566 528
rect 1520 446 1566 494
rect 1520 412 1526 446
rect 1560 412 1566 446
rect 1520 380 1566 412
rect 1630 596 2380 608
rect 1630 562 1636 596
rect 1670 562 1988 596
rect 2022 562 2340 596
rect 2374 562 2380 596
rect 1630 504 1676 562
rect 1630 470 1636 504
rect 1670 470 1676 504
rect 1630 413 1676 470
rect 1630 379 1636 413
rect 1670 379 1676 413
rect 1630 367 1676 379
rect 1806 516 1852 528
rect 1806 482 1812 516
rect 1846 482 1852 516
rect 1806 426 1852 482
rect 1806 392 1812 426
rect 1846 392 1852 426
rect 1806 337 1852 392
rect 992 303 998 337
rect 1032 303 1350 337
rect 1384 303 1812 337
rect 1846 303 1852 337
rect 992 291 1852 303
rect 1982 509 2028 562
rect 1982 475 1988 509
rect 2022 475 2028 509
rect 1982 423 2028 475
rect 1982 389 1988 423
rect 2022 389 2028 423
rect 2154 526 2206 532
rect 2154 462 2206 474
rect 2154 404 2164 410
rect 1982 337 2028 389
rect 1982 303 1988 337
rect 2022 303 2028 337
rect 1982 291 2028 303
rect 2158 392 2164 404
rect 2198 404 2206 410
rect 2334 509 2380 562
rect 2334 475 2340 509
rect 2374 475 2380 509
rect 2334 423 2380 475
rect 2198 392 2204 404
rect 2158 337 2204 392
rect 2158 303 2164 337
rect 2198 303 2204 337
rect 2158 291 2204 303
rect 2334 389 2340 423
rect 2374 389 2380 423
rect 2334 337 2380 389
rect 2334 303 2340 337
rect 2374 303 2380 337
rect 2334 291 2380 303
rect 2444 577 2450 611
rect 2484 577 2490 611
rect 2796 611 2842 643
rect 2444 526 2490 577
rect 2620 596 2666 608
rect 2620 562 2626 596
rect 2660 562 2666 596
rect 2444 492 2450 526
rect 2484 492 2490 526
rect 2444 441 2490 492
rect 2444 407 2450 441
rect 2484 407 2490 441
rect 2444 357 2490 407
rect 2539 526 2591 532
rect 2539 462 2591 474
rect 2539 404 2591 410
rect 2620 509 2666 562
rect 2620 475 2626 509
rect 2660 475 2666 509
rect 2620 423 2666 475
rect 2444 323 2450 357
rect 2484 323 2490 357
rect 2444 291 2490 323
rect 2620 389 2626 423
rect 2660 389 2666 423
rect 2620 343 2666 389
rect 2796 577 2802 611
rect 2836 577 2842 611
rect 3148 611 3194 643
rect 2796 528 2842 577
rect 2972 596 3018 608
rect 2972 570 2978 596
rect 3012 570 3018 596
rect 3148 577 3154 611
rect 3188 577 3194 611
rect 3500 611 3546 643
rect 2796 494 2802 528
rect 2836 494 2842 528
rect 2796 445 2842 494
rect 2796 411 2802 445
rect 2836 411 2842 445
rect 2796 379 2842 411
rect 2886 562 2978 570
rect 2886 518 2997 562
rect 3049 518 3061 570
rect 3113 518 3119 570
rect 2886 509 3119 518
rect 2886 475 2978 509
rect 3012 475 3119 509
rect 2886 423 3119 475
rect 2886 389 2978 423
rect 3012 389 3119 423
rect 2886 343 3119 389
rect 3148 528 3194 577
rect 3148 494 3154 528
rect 3188 494 3194 528
rect 3148 445 3194 494
rect 3148 411 3154 445
rect 3188 411 3194 445
rect 3148 379 3194 411
rect 3324 596 3370 608
rect 3324 562 3330 596
rect 3364 562 3370 596
rect 3324 509 3370 562
rect 3324 475 3330 509
rect 3364 475 3370 509
rect 3324 423 3370 475
rect 3324 389 3330 423
rect 3364 389 3370 423
rect 3324 343 3370 389
rect 2620 337 3370 343
rect 2620 303 2626 337
rect 2660 303 2978 337
rect 3012 303 3330 337
rect 3364 303 3370 337
rect 2620 291 3370 303
rect 3500 577 3506 611
rect 3540 577 3546 611
rect 3852 611 3898 643
rect 3500 521 3546 577
rect 3500 487 3506 521
rect 3540 487 3546 521
rect 3676 596 3722 608
rect 3676 562 3682 596
rect 3716 562 3722 596
rect 3676 518 3722 562
rect 3852 577 3858 611
rect 3892 577 3898 611
rect 4204 611 4250 643
rect 3852 528 3898 577
rect 3675 509 3803 518
rect 3675 506 3682 509
rect 3716 506 3803 509
rect 3500 431 3546 487
rect 3674 454 3680 506
rect 3732 454 3744 506
rect 3796 454 3803 506
rect 3500 397 3506 431
rect 3540 397 3546 431
rect 3500 341 3546 397
rect 3500 307 3506 341
rect 3540 307 3546 341
rect 3500 275 3546 307
rect 3675 423 3803 454
rect 3675 389 3682 423
rect 3716 389 3803 423
rect 3675 338 3803 389
rect 3852 494 3858 528
rect 3892 494 3898 528
rect 3852 445 3898 494
rect 3852 411 3858 445
rect 3892 411 3898 445
rect 3852 379 3898 411
rect 4028 596 4074 608
rect 4028 562 4034 596
rect 4068 562 4074 596
rect 4028 509 4074 562
rect 4028 475 4034 509
rect 4068 475 4074 509
rect 4028 423 4074 475
rect 4028 389 4034 423
rect 4068 389 4074 423
rect 4028 338 4074 389
rect 4204 577 4210 611
rect 4244 577 4250 611
rect 4908 611 4954 643
rect 4204 528 4250 577
rect 4204 494 4210 528
rect 4244 494 4250 528
rect 4204 445 4250 494
rect 4204 411 4210 445
rect 4244 411 4250 445
rect 4204 379 4250 411
rect 4380 596 4426 608
rect 4380 562 4386 596
rect 4420 562 4426 596
rect 4380 509 4426 562
rect 4380 475 4386 509
rect 4420 475 4426 509
rect 4732 596 4778 608
rect 4732 562 4738 596
rect 4772 562 4778 596
rect 4732 509 4778 562
rect 4380 423 4426 475
rect 4380 389 4386 423
rect 4420 389 4426 423
rect 4380 338 4426 389
rect 3675 337 4426 338
rect 3675 303 3682 337
rect 3716 303 4034 337
rect 4068 303 4386 337
rect 4420 303 4426 337
rect 3675 291 4426 303
rect 4566 453 4572 505
rect 4624 453 4636 505
rect 4688 453 4694 505
rect 4566 343 4694 453
rect 4732 475 4738 509
rect 4772 475 4778 509
rect 4732 423 4778 475
rect 4732 389 4738 423
rect 4772 389 4778 423
rect 4732 343 4778 389
rect 4908 577 4914 611
rect 4948 577 4954 611
rect 5260 611 5306 643
rect 4908 528 4954 577
rect 4908 494 4914 528
rect 4948 494 4954 528
rect 4908 445 4954 494
rect 4908 411 4914 445
rect 4948 411 4954 445
rect 4908 379 4954 411
rect 5084 596 5130 608
rect 5084 562 5090 596
rect 5124 562 5130 596
rect 5084 509 5130 562
rect 5084 475 5090 509
rect 5124 475 5130 509
rect 5084 423 5130 475
rect 5084 389 5090 423
rect 5124 389 5130 423
rect 5084 343 5130 389
rect 5260 577 5266 611
rect 5300 577 5306 611
rect 5612 611 5658 643
rect 5260 528 5306 577
rect 5260 494 5266 528
rect 5300 494 5306 528
rect 5260 445 5306 494
rect 5260 411 5266 445
rect 5300 411 5306 445
rect 5260 379 5306 411
rect 5436 596 5482 608
rect 5436 562 5442 596
rect 5476 562 5482 596
rect 5436 509 5482 562
rect 5436 475 5442 509
rect 5476 475 5482 509
rect 5436 423 5482 475
rect 5436 389 5442 423
rect 5476 389 5482 423
rect 5436 343 5482 389
rect 5612 577 5618 611
rect 5652 577 5658 611
rect 5612 521 5658 577
rect 5612 487 5618 521
rect 5652 487 5658 521
rect 5612 431 5658 487
rect 5612 397 5618 431
rect 5652 397 5658 431
rect 4566 337 5526 343
rect 4566 303 4738 337
rect 4772 303 5090 337
rect 5124 303 5442 337
rect 5476 303 5526 337
rect 4566 291 5526 303
rect 5612 341 5658 397
rect 5612 307 5618 341
rect 5652 307 5658 341
rect 3675 286 4425 291
rect 5612 275 5658 307
<< via1 >>
rect 266 1882 382 1998
rect 2539 1613 2591 1665
rect 2539 1549 2591 1601
rect 2997 1507 3049 1559
rect 3061 1556 3113 1559
rect 3061 1522 3097 1556
rect 3097 1522 3113 1556
rect 3061 1507 3113 1522
rect 1169 1432 1221 1484
rect 1233 1432 1285 1484
rect 2823 1425 2875 1477
rect 2887 1425 2939 1477
rect 4572 1425 4624 1477
rect 4636 1425 4688 1477
rect 6122 1317 6174 1357
rect 6122 1305 6134 1317
rect 6134 1305 6168 1317
rect 6168 1305 6174 1317
rect 6122 1235 6174 1247
rect 6122 1201 6134 1235
rect 6134 1201 6168 1235
rect 6168 1201 6174 1235
rect 6122 1195 6174 1201
rect 1163 1145 1215 1151
rect 1163 1111 1175 1145
rect 1175 1111 1209 1145
rect 1209 1111 1215 1145
rect 1163 1099 1215 1111
rect 2124 1142 2176 1148
rect 2188 1142 2240 1148
rect 2124 1108 2137 1142
rect 2137 1108 2175 1142
rect 2175 1108 2176 1142
rect 2188 1108 2209 1142
rect 2209 1108 2240 1142
rect 2124 1096 2176 1108
rect 2188 1096 2240 1108
rect 2823 1142 2875 1148
rect 2823 1108 2853 1142
rect 2853 1108 2875 1142
rect 2823 1096 2875 1108
rect 2887 1142 2939 1148
rect 2887 1108 2891 1142
rect 2891 1108 2925 1142
rect 2925 1108 2939 1142
rect 2887 1096 2939 1108
rect 4982 1142 5034 1148
rect 4982 1108 5009 1142
rect 5009 1108 5034 1142
rect 4982 1096 5034 1108
rect 5046 1142 5098 1148
rect 5046 1108 5047 1142
rect 5047 1108 5081 1142
rect 5081 1108 5098 1142
rect 5046 1096 5098 1108
rect 1163 1073 1215 1087
rect 1163 1039 1175 1073
rect 1175 1039 1209 1073
rect 1209 1039 1215 1073
rect 1163 1035 1215 1039
rect 1163 971 1215 1023
rect 5770 1062 5822 1068
rect 5880 1062 5932 1068
rect 5770 1028 5807 1062
rect 5807 1028 5822 1062
rect 5880 1028 5913 1062
rect 5913 1028 5932 1062
rect 5770 1016 5822 1028
rect 5880 1016 5932 1028
rect 2346 915 2398 967
rect 2410 915 2462 967
rect 4393 915 4445 967
rect 4457 915 4509 967
rect 4982 961 5034 967
rect 4982 927 5012 961
rect 5012 927 5034 961
rect 4982 915 5034 927
rect 5046 961 5098 967
rect 5046 927 5050 961
rect 5050 927 5084 961
rect 5084 927 5098 961
rect 5046 915 5098 927
rect 266 799 360 833
rect 360 799 382 833
rect 266 761 382 799
rect 266 727 360 761
rect 360 727 382 761
rect 266 689 382 727
rect 266 655 360 689
rect 360 655 382 689
rect 266 653 382 655
rect 266 478 382 594
rect 2154 516 2206 526
rect 2154 482 2164 516
rect 2164 482 2198 516
rect 2198 482 2206 516
rect 2154 474 2206 482
rect 2154 426 2206 462
rect 2154 410 2164 426
rect 2164 410 2198 426
rect 2198 410 2206 426
rect 2539 474 2591 526
rect 2539 410 2591 462
rect 2997 562 3012 570
rect 3012 562 3049 570
rect 2997 518 3049 562
rect 3061 518 3113 570
rect 3680 475 3682 506
rect 3682 475 3716 506
rect 3716 475 3732 506
rect 3680 454 3732 475
rect 3744 454 3796 506
rect 4572 453 4624 505
rect 4636 453 4688 505
<< metal2 >>
rect 260 1998 388 2005
rect 260 1882 266 1998
rect 382 1882 388 1998
rect 260 833 388 1882
rect 2539 1665 2591 1692
rect 2539 1601 2591 1613
rect 1163 1432 1169 1484
rect 1221 1432 1233 1484
rect 1285 1432 1291 1484
rect 1163 1425 1233 1432
tri 1233 1425 1240 1432 nw
rect 1163 1151 1215 1425
tri 1215 1407 1233 1425 nw
rect 1163 1087 1215 1099
rect 1163 1023 1215 1035
rect 1163 965 1215 971
rect 2118 1096 2124 1148
rect 2176 1096 2188 1148
rect 2240 1096 2246 1148
rect 2118 974 2246 1096
rect 2118 967 2468 974
rect 260 653 266 833
rect 382 653 388 833
rect 260 594 388 653
rect 260 478 266 594
rect 382 478 388 594
rect 2118 915 2346 967
rect 2398 915 2410 967
rect 2462 915 2468 967
rect 2118 913 2468 915
rect 2118 526 2207 913
tri 2207 874 2246 913 nw
rect 2118 474 2154 526
rect 2206 474 2207 526
rect 2118 462 2207 474
rect 2118 410 2154 462
rect 2206 410 2207 462
rect 2118 404 2207 410
rect 2539 526 2591 1549
rect 2991 1507 2997 1559
rect 3049 1507 3061 1559
rect 3113 1507 3119 1559
rect 2817 1425 2823 1477
rect 2875 1425 2887 1477
rect 2939 1425 2945 1477
rect 2817 1148 2945 1425
rect 2817 1096 2823 1148
rect 2875 1096 2887 1148
rect 2939 1096 2945 1148
rect 2991 570 3119 1507
rect 4566 1425 4572 1477
rect 4624 1425 4636 1477
rect 4688 1425 4694 1477
rect 2991 518 2997 570
rect 3049 518 3061 570
rect 3113 518 3119 570
rect 4387 915 4393 967
rect 4445 915 4457 967
rect 4509 915 4515 967
rect 3674 488 3680 506
rect 2591 474 3680 488
rect 2539 462 3680 474
rect 2591 454 3680 462
rect 3732 454 3744 506
rect 3796 488 3802 506
rect 4387 488 4515 915
rect 3796 454 4515 488
rect 4566 505 4694 1425
tri 5820 1357 5826 1363 se
rect 5826 1357 6174 1363
tri 5768 1305 5820 1357 se
rect 5820 1305 6122 1357
tri 5764 1301 5768 1305 se
rect 5768 1301 6174 1305
rect 5764 1247 6174 1301
rect 5764 1195 6122 1247
rect 5764 1189 6174 1195
rect 4976 1096 4982 1148
rect 5034 1096 5046 1148
rect 5098 1096 5104 1148
rect 4976 967 5104 1096
rect 5764 1068 5938 1189
rect 5764 1016 5770 1068
rect 5822 1016 5880 1068
rect 5932 1016 5938 1068
rect 4976 915 4982 967
rect 5034 915 5046 967
rect 5098 915 5104 967
rect 4566 453 4572 505
rect 4624 453 4636 505
rect 4688 453 4694 505
rect 2539 404 2591 410
use sky130_fd_pr__nfet_01v8__example_55959141808360  sky130_fd_pr__nfet_01v8__example_55959141808360_0
timestamp 1679235063
transform -1 0 811 0 1 279
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808362  sky130_fd_pr__nfet_01v8__example_55959141808362_0
timestamp 1679235063
transform 1 0 2033 0 1 279
box -1 0 297 1
use sky130_fd_pr__nfet_01v8__example_55959141808362  sky130_fd_pr__nfet_01v8__example_55959141808362_1
timestamp 1679235063
transform 1 0 1681 0 1 279
box -1 0 297 1
use sky130_fd_pr__nfet_01v8__example_55959141808403  sky130_fd_pr__nfet_01v8__example_55959141808403_0
timestamp 1679235063
transform -1 0 1515 0 1 279
box -1 0 649 1
use sky130_fd_pr__nfet_01v8__example_55959141808404  sky130_fd_pr__nfet_01v8__example_55959141808404_0
timestamp 1679235063
transform -1 0 3495 0 1 279
box -1 0 1001 1
use sky130_fd_pr__nfet_01v8__example_55959141808404  sky130_fd_pr__nfet_01v8__example_55959141808404_1
timestamp 1679235063
transform 1 0 3551 0 1 279
box -1 0 1001 1
use sky130_fd_pr__nfet_01v8__example_55959141808405  sky130_fd_pr__nfet_01v8__example_55959141808405_0
timestamp 1679235063
transform 1 0 405 0 1 279
box -1 0 121 1
use sky130_fd_pr__nfet_01v8__example_55959141808406  sky130_fd_pr__nfet_01v8__example_55959141808406_0
timestamp 1679235063
transform 1 0 4607 0 1 279
box -1 0 297 1
use sky130_fd_pr__nfet_01v8__example_55959141808406  sky130_fd_pr__nfet_01v8__example_55959141808406_1
timestamp 1679235063
transform 1 0 5311 0 1 279
box -1 0 297 1
use sky130_fd_pr__nfet_01v8__example_55959141808406  sky130_fd_pr__nfet_01v8__example_55959141808406_2
timestamp 1679235063
transform 1 0 4959 0 1 279
box -1 0 297 1
use sky130_fd_pr__pfet_01v8__example_55959141808346  sky130_fd_pr__pfet_01v8__example_55959141808346_0
timestamp 1679235063
transform -1 0 6007 0 -1 2193
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808346  sky130_fd_pr__pfet_01v8__example_55959141808346_1
timestamp 1679235063
transform 1 0 4815 0 -1 2193
box -1 0 569 1
use sky130_fd_pr__pfet_01v8__example_55959141808407  sky130_fd_pr__pfet_01v8__example_55959141808407_0
timestamp 1679235063
transform -1 0 3241 0 -1 2193
box -1 0 881 1
use sky130_fd_pr__pfet_01v8__example_55959141808408  sky130_fd_pr__pfet_01v8__example_55959141808408_0
timestamp 1679235063
transform 1 0 3297 0 -1 2193
box -1 0 1353 1
use sky130_fd_pr__pfet_01v8__example_55959141808409  sky130_fd_pr__pfet_01v8__example_55959141808409_0
timestamp 1679235063
transform 1 0 691 0 -1 2193
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808409  sky130_fd_pr__pfet_01v8__example_55959141808409_1
timestamp 1679235063
transform -1 0 947 0 -1 2193
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808409  sky130_fd_pr__pfet_01v8__example_55959141808409_2
timestamp 1679235063
transform 1 0 1159 0 -1 2193
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808409  sky130_fd_pr__pfet_01v8__example_55959141808409_3
timestamp 1679235063
transform -1 0 1103 0 -1 2193
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808409  sky130_fd_pr__pfet_01v8__example_55959141808409_4
timestamp 1679235063
transform 1 0 405 0 -1 2193
box -1 0 101 1
use sky130_fd_pr__pfet_01v8__example_55959141808410  sky130_fd_pr__pfet_01v8__example_55959141808410_0
timestamp 1679235063
transform -1 0 2305 0 -1 2193
box -1 0 881 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1679235063
transform 0 -1 924 -1 0 1145
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1679235063
transform -1 0 570 0 1 1194
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1679235063
transform 0 -1 1070 -1 0 1145
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1679235063
transform 1 0 622 0 1 879
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1679235063
transform 0 -1 1209 -1 0 1145
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1679235063
transform 0 -1 5300 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1679235063
transform 0 -1 5652 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_2
timestamp 1679235063
transform 0 -1 4948 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_3
timestamp 1679235063
transform 0 -1 4596 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_4
timestamp 1679235063
transform 0 -1 4244 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_5
timestamp 1679235063
transform 0 -1 3892 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_6
timestamp 1679235063
transform 0 -1 3540 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_7
timestamp 1679235063
transform 0 -1 3188 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_8
timestamp 1679235063
transform 0 -1 2836 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_9
timestamp 1679235063
transform 0 -1 2484 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_10
timestamp 1679235063
transform 0 -1 856 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_11
timestamp 1679235063
transform 0 -1 1208 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_12
timestamp 1679235063
transform 0 -1 1560 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_13
timestamp 1679235063
transform 0 -1 6168 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_14
timestamp 1679235063
transform 0 -1 394 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_15
timestamp 1679235063
transform 0 -1 394 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_16
timestamp 1679235063
transform 0 -1 836 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_17
timestamp 1679235063
transform 0 -1 1148 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_18
timestamp 1679235063
transform 0 -1 1414 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_19
timestamp 1679235063
transform 0 -1 1726 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_20
timestamp 1679235063
transform 0 -1 2038 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_21
timestamp 1679235063
transform 0 -1 2350 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_22
timestamp 1679235063
transform 0 -1 3638 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_23
timestamp 1679235063
transform 0 -1 3286 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_24
timestamp 1679235063
transform 0 -1 2974 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_25
timestamp 1679235063
transform 0 -1 2662 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_26
timestamp 1679235063
transform 0 -1 3990 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_27
timestamp 1679235063
transform 0 -1 4342 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_28
timestamp 1679235063
transform 0 -1 4694 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_29
timestamp 1679235063
transform 0 -1 5768 1 0 655
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_30
timestamp 1679235063
transform 0 -1 122 1 0 2045
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_0
timestamp 1679235063
transform 1 0 196 0 1 1120
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_1
timestamp 1679235063
transform -1 0 5228 0 1 927
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_2
timestamp 1679235063
transform -1 0 1955 0 1 954
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808127  sky130_fd_pr__via_l1m1__example_55959141808127_3
timestamp 1679235063
transform -1 0 2298 0 1 879
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808269  sky130_fd_pr__via_l1m1__example_55959141808269_0
timestamp 1679235063
transform 1 0 3350 0 1 1108
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808290  sky130_fd_pr__via_l1m1__example_55959141808290_0
timestamp 1679235063
transform 1 0 4831 0 1 1108
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808325  sky130_fd_pr__via_l1m1__example_55959141808325_0
timestamp 1679235063
transform 1 0 1289 0 1 1028
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808326  sky130_fd_pr__via_l1m1__example_55959141808326_0
timestamp 1679235063
transform -1 0 4317 0 1 927
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808372  sky130_fd_pr__via_l1m1__example_55959141808372_0
timestamp 1679235063
transform 1 0 5663 0 1 1028
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808399  sky130_fd_pr__via_l1m1__example_55959141808399_0
timestamp 1679235063
transform 1 0 3298 0 1 1028
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808400  sky130_fd_pr__via_l1m1__example_55959141808400_0
timestamp 1679235063
transform 1 0 1455 0 1 1108
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808400  sky130_fd_pr__via_l1m1__example_55959141808400_1
timestamp 1679235063
transform -1 0 3213 0 1 1108
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_55959141808401  sky130_fd_pr__via_l1m1__example_55959141808401_0
timestamp 1679235063
transform 1 0 -99 0 1 484
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_0
timestamp 1679235063
transform 0 -1 2591 1 0 404
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_1
timestamp 1679235063
transform 0 -1 2206 1 0 404
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_2
timestamp 1679235063
transform 1 0 2340 0 -1 967
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_3
timestamp 1679235063
transform 1 0 2991 0 1 518
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_4
timestamp 1679235063
transform 1 0 2991 0 1 1507
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_5
timestamp 1679235063
transform 1 0 1163 0 1 1432
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_6
timestamp 1679235063
transform 1 0 3674 0 1 454
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_7
timestamp 1679235063
transform 1 0 2118 0 -1 1148
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_8
timestamp 1679235063
transform -1 0 4515 0 1 915
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_9
timestamp 1679235063
transform -1 0 5104 0 1 915
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_10
timestamp 1679235063
transform -1 0 5104 0 1 1096
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_11
timestamp 1679235063
transform 1 0 4566 0 1 1425
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_12
timestamp 1679235063
transform 1 0 4566 0 1 453
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_13
timestamp 1679235063
transform -1 0 2945 0 1 1425
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808260  sky130_fd_pr__via_m1m2__example_55959141808260_14
timestamp 1679235063
transform -1 0 2945 0 -1 1148
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808261  sky130_fd_pr__via_m1m2__example_55959141808261_0
timestamp 1679235063
transform 0 -1 1215 -1 0 1157
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_0
timestamp 1679235063
transform 1 0 260 0 1 1882
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808350  sky130_fd_pr__via_m1m2__example_55959141808350_1
timestamp 1679235063
transform 1 0 260 0 1 478
box 0 0 1 1
use sky130_fd_pr__via_m1m2__example_55959141808402  sky130_fd_pr__via_m1m2__example_55959141808402_0
timestamp 1679235063
transform 1 0 260 0 1 653
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_0
timestamp 1679235063
transform 1 0 1020 0 1 1027
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_1
timestamp 1679235063
transform 1 0 874 0 -1 1145
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_2
timestamp 1679235063
transform 1 0 1159 0 -1 1161
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_5595914180833  sky130_fd_pr__via_pol1__example_5595914180833_3
timestamp 1679235063
transform 1 0 704 0 -1 1145
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808274  sky130_fd_pr__via_pol1__example_55959141808274_0
timestamp 1679235063
transform -1 0 486 0 -1 1158
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_0
timestamp 1679235063
transform 0 1 5455 -1 0 1161
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808294  sky130_fd_pr__via_pol1__example_55959141808294_1
timestamp 1679235063
transform 0 1 4819 -1 0 1161
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808295  sky130_fd_pr__via_pol1__example_55959141808295_0
timestamp 1679235063
transform 0 1 884 -1 0 985
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_0
timestamp 1679235063
transform 0 -1 2318 -1 0 977
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_1
timestamp 1679235063
transform 0 -1 1971 -1 0 977
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808298  sky130_fd_pr__via_pol1__example_55959141808298_2
timestamp 1679235063
transform 0 1 5322 1 0 911
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808322  sky130_fd_pr__via_pol1__example_55959141808322_0
timestamp 1679235063
transform 0 -1 2281 -1 0 1161
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808322  sky130_fd_pr__via_pol1__example_55959141808322_1
timestamp 1679235063
transform 0 -1 3217 -1 0 1161
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808394  sky130_fd_pr__via_pol1__example_55959141808394_0
timestamp 1679235063
transform 0 -1 4529 -1 0 977
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808394  sky130_fd_pr__via_pol1__example_55959141808394_1
timestamp 1679235063
transform 0 -1 3479 -1 0 977
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808395  sky130_fd_pr__via_pol1__example_55959141808395_0
timestamp 1679235063
transform 1 0 5439 0 1 1027
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808396  sky130_fd_pr__via_pol1__example_55959141808396_0
timestamp 1679235063
transform 0 1 4970 1 0 911
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808396  sky130_fd_pr__via_pol1__example_55959141808396_1
timestamp 1679235063
transform 0 1 4618 1 0 911
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808397  sky130_fd_pr__via_pol1__example_55959141808397_0
timestamp 1679235063
transform 0 1 3319 -1 0 1161
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_55959141808398  sky130_fd_pr__via_pol1__example_55959141808398_0
timestamp 1679235063
transform -1 0 3241 0 1 1007
box 0 0 1 1
<< labels >>
flabel locali s 720 1111 754 1145 3 FreeSans 300 0 0 0 PU_DIS_H
port 1 nsew
flabel locali s 5947 1111 5997 1145 3 FreeSans 300 0 0 0 PD_DIS_H
port 2 nsew
flabel metal1 s 22 1875 62 2005 3 FreeSans 300 0 0 0 VGND
port 3 nsew
flabel metal1 s 303 1114 349 1160 3 FreeSans 300 0 0 0 OE_H
port 4 nsew
flabel metal1 s 1486 1543 1536 1595 3 FreeSans 300 180 0 0 DRVHI_H
port 6 nsew
flabel metal1 s 6229 648 6269 1156 3 FreeSans 300 180 0 0 VGND
port 3 nsew
flabel metal1 s 6194 2033 6234 2235 3 FreeSans 300 180 0 0 VCC_IO
port 7 nsew
flabel metal1 s -47 884 -7 1086 3 FreeSans 300 180 0 0 VGND
port 3 nsew
flabel metal1 s 22 2033 62 2235 3 FreeSans 300 180 0 0 VCC_IO
port 7 nsew
flabel metal1 s 6103 800 6143 930 3 FreeSans 300 180 0 0 VGND
port 3 nsew
flabel metal1 s 1163 1432 1215 1484 3 FreeSans 300 180 0 0 DRVLO_H_N
port 5 nsew
flabel metal1 s 1189 1458 1189 1458 3 FreeSans 300 180 0 0 DRVLO_H_N
flabel comment s 5095 971 5095 971 0 FreeSans 300 0 0 0 DRVHI_H
flabel comment s 4861 593 4861 593 0 FreeSans 300 180 0 0 N1
flabel comment s 31 2217 31 2217 0 FreeSans 300 0 0 0 VCC_IO
flabel comment s 1696 1748 1696 1748 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 2486 1748 2486 1748 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 4387 1828 4387 1828 0 FreeSans 300 0 0 0 DRVHI_H
flabel comment s 3050 1828 3050 1828 0 FreeSans 300 0 0 0 DRVHI_H
flabel comment s 4722 1065 4722 1065 0 FreeSans 300 180 0 0 OE_I_H_N
flabel comment s 4157 1756 4157 1756 0 FreeSans 300 180 0 0 INT_NOR_N<0>
flabel comment s 4906 1825 4906 1825 0 FreeSans 300 180 0 0 INT_NOR_N<1>
flabel comment s 1233 1663 1233 1663 0 FreeSans 300 180 0 0 N0
flabel comment s 2238 596 2238 596 0 FreeSans 300 0 0 0 N0
flabel comment s 1712 509 1712 509 0 FreeSans 300 0 0 0 INT_NAND_N1
flabel comment s 1069 600 1069 600 0 FreeSans 300 0 0 0 INT_NAND_N0
flabel comment s 3108 1748 3108 1748 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 5673 1665 5673 1665 0 FreeSans 300 180 0 0 N1
flabel comment s 2777 505 2777 505 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 3833 505 3833 505 0 FreeSans 300 0 0 0 DRVHI_H
flabel comment s 2946 986 2946 986 0 FreeSans 300 180 0 0 N1
flabel comment s 740 904 740 904 0 FreeSans 300 270 0 0 PU_DIS_H
flabel comment s 1823 984 1823 984 0 FreeSans 300 0 0 0 DRVLO_H_N
flabel comment s 1161 984 1161 984 0 FreeSans 300 0 0 0 OE_I_H
flabel comment s 3804 977 3804 977 0 FreeSans 300 180 0 0 N0
flabel comment s 5446 975 5446 975 0 FreeSans 300 180 0 0 PD_DIS_H
flabel comment s 1808 1828 1808 1828 0 FreeSans 300 0 0 0 DRVHI_H
flabel comment s 2214 986 2214 986 0 FreeSans 300 0 0 0 PU_DIS_H_N
flabel comment s 536 1006 536 1006 0 FreeSans 300 90 0 0 OE_I_H_N
flabel comment s 4016 1098 4016 1098 0 FreeSans 300 180 0 0 OE_I_H_N
flabel comment s 4863 1097 4863 1097 0 FreeSans 300 180 0 0 DRVHI_H
flabel comment s 2803 1098 2803 1098 0 FreeSans 300 180 0 0 N1
flabel comment s 1024 1139 1024 1139 0 FreeSans 300 90 0 0 PU_DIS_H_N
flabel comment s 1851 1155 1851 1155 0 FreeSans 300 180 0 0 N0
flabel comment s 1165 1134 1165 1134 0 FreeSans 300 90 0 0 DRVLO_H_N
flabel comment s 892 920 892 920 0 FreeSans 300 90 0 0 OE_I_H
flabel comment s 449 898 449 898 0 FreeSans 300 90 0 0 OE_I_H
flabel comment s 5733 1093 5733 1093 0 FreeSans 300 180 0 0 PD_DIS_H
<< properties >>
string GDS_END 36803084
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 36737412
<< end >>
