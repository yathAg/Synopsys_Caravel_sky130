magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1173 157 1355 201
rect 1661 157 2390 203
rect 1 145 825 157
rect 1027 145 2390 157
rect 1 21 2390 145
rect 29 -17 63 21
<< locali >>
rect 19 195 89 325
rect 356 157 390 337
rect 492 271 559 337
rect 617 157 651 223
rect 707 207 807 331
rect 356 123 651 157
rect 495 61 530 123
rect 1851 306 1917 486
rect 1851 299 1923 306
rect 1882 286 1923 299
rect 1889 178 1923 286
rect 1882 165 1923 178
rect 1851 158 1923 165
rect 2238 289 2288 465
rect 1851 51 1917 158
rect 2247 159 2288 289
rect 2238 53 2288 159
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 36 393 70 493
rect 104 427 170 527
rect 36 359 169 393
rect 123 194 169 359
rect 123 161 162 194
rect 35 127 162 161
rect 204 143 249 493
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 249 143
rect 287 415 342 489
rect 376 449 442 527
rect 539 449 718 483
rect 287 372 650 415
rect 287 89 321 372
rect 424 225 458 372
rect 616 337 650 372
rect 684 399 718 449
rect 752 433 786 527
rect 841 413 897 488
rect 937 438 1151 472
rect 841 399 875 413
rect 684 365 875 399
rect 616 271 655 337
rect 424 191 493 225
rect 841 173 875 365
rect 685 139 875 173
rect 909 207 957 381
rect 995 331 1083 402
rect 1117 315 1151 438
rect 1185 367 1219 527
rect 1253 427 1303 493
rect 1348 433 1525 467
rect 1117 297 1219 315
rect 1059 263 1219 297
rect 909 141 1025 207
rect 287 55 361 89
rect 395 17 461 89
rect 685 89 719 139
rect 841 107 875 139
rect 1059 107 1093 263
rect 1185 249 1219 263
rect 1127 213 1161 219
rect 1253 213 1287 427
rect 1321 249 1359 393
rect 1393 315 1457 381
rect 1127 153 1287 213
rect 1393 207 1431 315
rect 1491 281 1525 433
rect 1561 427 1622 527
rect 1679 381 1745 491
rect 1559 315 1745 381
rect 1779 325 1815 527
rect 564 55 719 89
rect 753 17 793 105
rect 841 73 911 107
rect 945 73 1093 107
rect 1143 17 1217 117
rect 1253 107 1287 153
rect 1321 141 1431 207
rect 1465 265 1525 281
rect 1708 265 1745 315
rect 1953 323 1987 527
rect 1465 199 1674 265
rect 1708 199 1855 265
rect 1465 107 1499 199
rect 1708 165 1745 199
rect 1253 73 1345 107
rect 1391 73 1499 107
rect 1548 17 1622 123
rect 1672 60 1745 165
rect 2041 265 2107 485
rect 2143 299 2204 527
rect 2041 199 2213 265
rect 1779 17 1817 139
rect 1951 17 1997 138
rect 2041 69 2091 199
rect 2138 17 2204 161
rect 2322 279 2356 527
rect 2322 17 2356 191
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< obsm1 >>
rect 117 388 175 397
rect 1029 388 1087 397
rect 1313 388 1371 397
rect 117 360 1371 388
rect 117 351 175 360
rect 1029 351 1087 360
rect 1313 351 1371 360
rect 198 184 256 193
rect 937 184 995 193
rect 1316 184 1374 193
rect 198 156 1374 184
rect 198 147 256 156
rect 937 147 995 156
rect 1316 147 1374 156
<< labels >>
rlabel locali s 19 195 89 325 6 CLK
port 1 nsew clock input
rlabel locali s 492 271 559 337 6 D
port 2 nsew signal input
rlabel locali s 707 207 807 331 6 SCD
port 3 nsew signal input
rlabel locali s 495 61 530 123 6 SCE
port 4 nsew signal input
rlabel locali s 356 123 651 157 6 SCE
port 4 nsew signal input
rlabel locali s 617 157 651 223 6 SCE
port 4 nsew signal input
rlabel locali s 356 157 390 337 6 SCE
port 4 nsew signal input
rlabel metal1 s 0 -48 2392 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 2390 145 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1027 145 2390 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 145 825 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1661 157 2390 203 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1173 157 1355 201 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 2430 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 2392 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1851 51 1917 158 6 Q
port 9 nsew signal output
rlabel locali s 1851 158 1923 165 6 Q
port 9 nsew signal output
rlabel locali s 1882 165 1923 178 6 Q
port 9 nsew signal output
rlabel locali s 1889 178 1923 286 6 Q
port 9 nsew signal output
rlabel locali s 1882 286 1923 299 6 Q
port 9 nsew signal output
rlabel locali s 1851 299 1923 306 6 Q
port 9 nsew signal output
rlabel locali s 1851 306 1917 486 6 Q
port 9 nsew signal output
rlabel locali s 2238 53 2288 159 6 Q_N
port 10 nsew signal output
rlabel locali s 2247 159 2288 289 6 Q_N
port 10 nsew signal output
rlabel locali s 2238 289 2288 465 6 Q_N
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2392 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 361040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 343158
<< end >>
