magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< locali >>
rect 12028 18138 12590 18733
rect 1835 1730 2397 2325
rect 1835 -41064 2397 -40469
<< obsli1 >>
rect 17363 20659 17497 20675
rect 17363 20625 17377 20659
rect 17411 20625 17449 20659
rect 17483 20625 17497 20659
rect 17363 20609 17497 20625
rect 18079 20659 18349 20675
rect 18079 20625 18089 20659
rect 18123 20625 18161 20659
rect 18195 20625 18233 20659
rect 18267 20625 18305 20659
rect 18339 20625 18349 20659
rect 18079 20609 18349 20625
rect 18915 20659 19457 20675
rect 18915 20625 18917 20659
rect 18951 20625 18989 20659
rect 19023 20625 19061 20659
rect 19095 20625 19133 20659
rect 19167 20625 19205 20659
rect 19239 20625 19277 20659
rect 19311 20625 19349 20659
rect 19383 20625 19421 20659
rect 19455 20625 19457 20659
rect 18915 20609 19457 20625
rect 17327 20547 17361 20563
rect 17327 20475 17361 20513
rect 17327 20403 17361 20441
rect 17327 20331 17361 20369
rect 17327 20259 17361 20297
rect 14875 20227 15009 20243
rect 14875 20193 14889 20227
rect 14923 20193 14961 20227
rect 14995 20193 15009 20227
rect 14875 20177 15009 20193
rect 15437 20227 15707 20243
rect 15437 20193 15447 20227
rect 15481 20193 15519 20227
rect 15553 20193 15591 20227
rect 15625 20193 15663 20227
rect 15697 20193 15707 20227
rect 15437 20177 15707 20193
rect 16116 20227 16658 20243
rect 16116 20193 16118 20227
rect 16152 20193 16190 20227
rect 16224 20193 16262 20227
rect 16296 20193 16334 20227
rect 16368 20193 16406 20227
rect 16440 20193 16478 20227
rect 16512 20193 16550 20227
rect 16584 20193 16622 20227
rect 16656 20193 16658 20227
rect 16116 20177 16658 20193
rect 17327 20187 17361 20225
rect 13851 20143 13985 20159
rect 13851 20109 13865 20143
rect 13899 20109 13937 20143
rect 13971 20109 13985 20143
rect 13851 20093 13985 20109
rect 14839 20115 14873 20131
rect 13815 20043 13849 20059
rect 13815 19993 13849 20009
rect 13901 19993 13935 20059
rect 13987 20043 14021 20059
rect 13987 19993 14021 20009
rect 14839 20043 14873 20081
rect 14839 19993 14873 20009
rect 14925 19993 14959 20131
rect 15011 20115 15045 20131
rect 15011 20043 15045 20081
rect 15011 19993 15045 20009
rect 15383 20115 15417 20131
rect 15383 20043 15417 20081
rect 15383 19993 15417 20009
rect 15469 19993 15503 20131
rect 15555 20115 15589 20131
rect 15555 20043 15589 20081
rect 15555 19993 15589 20009
rect 15641 19993 15675 20131
rect 15727 20115 15761 20131
rect 15727 20043 15761 20081
rect 15727 19993 15761 20009
rect 16026 20115 16060 20131
rect 16026 20043 16060 20081
rect 16026 19993 16060 20009
rect 16112 19993 16146 20131
rect 16198 20115 16232 20131
rect 16198 20043 16232 20081
rect 16198 19993 16232 20009
rect 16284 19993 16318 20131
rect 16370 20115 16404 20131
rect 16370 20043 16404 20081
rect 16370 19993 16404 20009
rect 16456 19993 16490 20131
rect 16542 20115 16576 20131
rect 16542 20043 16576 20081
rect 16542 19993 16576 20009
rect 16628 19993 16662 20131
rect 16714 20115 16748 20131
rect 16714 20043 16748 20081
rect 16714 19993 16748 20009
rect 17327 20115 17361 20153
rect 17327 20043 17361 20081
rect 17327 19989 17361 20009
rect 17413 19993 17447 20563
rect 17499 20547 17533 20563
rect 17499 20475 17533 20513
rect 17499 20403 17533 20441
rect 17499 20331 17533 20369
rect 17499 20259 17533 20297
rect 17499 20187 17533 20225
rect 17499 20115 17533 20153
rect 17499 20043 17533 20081
rect 17499 19993 17533 20009
rect 18025 20547 18059 20563
rect 18025 20475 18059 20513
rect 18025 20403 18059 20441
rect 18025 20331 18059 20369
rect 18025 20259 18059 20297
rect 18025 20187 18059 20225
rect 18025 20115 18059 20153
rect 18025 20043 18059 20081
rect 18025 19993 18059 20009
rect 18111 19993 18145 20563
rect 18197 20547 18231 20563
rect 18197 20475 18231 20513
rect 18197 20403 18231 20441
rect 18197 20331 18231 20369
rect 18197 20259 18231 20297
rect 18197 20187 18231 20225
rect 18197 20115 18231 20153
rect 18197 20043 18231 20081
rect 18197 19993 18231 20009
rect 18283 19993 18317 20563
rect 18369 20547 18403 20563
rect 18369 20475 18403 20513
rect 18369 20403 18403 20441
rect 18369 20331 18403 20369
rect 18369 20259 18403 20297
rect 18369 20187 18403 20225
rect 18369 20115 18403 20153
rect 18369 20043 18403 20081
rect 18369 19993 18403 20009
rect 18825 20547 18859 20563
rect 18825 20475 18859 20513
rect 18825 20403 18859 20441
rect 18825 20331 18859 20369
rect 18825 20259 18859 20297
rect 18825 20187 18859 20225
rect 18825 20115 18859 20153
rect 18825 20043 18859 20081
rect 18825 19993 18859 20009
rect 18911 19993 18945 20563
rect 18997 20547 19031 20563
rect 18997 20475 19031 20513
rect 18997 20403 19031 20441
rect 18997 20331 19031 20369
rect 18997 20259 19031 20297
rect 18997 20187 19031 20225
rect 18997 20115 19031 20153
rect 18997 20043 19031 20081
rect 18997 19993 19031 20009
rect 19083 19993 19117 20563
rect 19169 20547 19203 20563
rect 19169 20475 19203 20513
rect 19169 20403 19203 20441
rect 19169 20331 19203 20369
rect 19169 20259 19203 20297
rect 19169 20187 19203 20225
rect 19169 20115 19203 20153
rect 19169 20043 19203 20081
rect 19169 19993 19203 20009
rect 19255 19993 19289 20563
rect 19341 20547 19375 20563
rect 19341 20475 19375 20513
rect 19341 20403 19375 20441
rect 19341 20331 19375 20369
rect 19341 20259 19375 20297
rect 19341 20187 19375 20225
rect 19341 20115 19375 20153
rect 19341 20043 19375 20081
rect 19341 19993 19375 20009
rect 19427 19993 19461 20563
rect 19513 20547 19547 20563
rect 19513 20475 19547 20513
rect 19513 20403 19547 20441
rect 19513 20331 19547 20369
rect 19513 20259 19547 20297
rect 19513 20187 19547 20225
rect 19513 20115 19547 20153
rect 19513 20043 19547 20081
rect 19513 19993 19547 20009
rect 17315 -23976 17449 -23960
rect 17315 -24010 17329 -23976
rect 17363 -24010 17401 -23976
rect 17435 -24010 17449 -23976
rect 17315 -24026 17449 -24010
rect 17279 -24109 17313 -24060
rect 17279 -24181 17313 -24143
rect 17279 -24253 17313 -24215
rect 17279 -24325 17313 -24287
rect 16432 -24383 16566 -24367
rect 16432 -24417 16446 -24383
rect 16480 -24417 16518 -24383
rect 16552 -24417 16566 -24383
rect 16432 -24435 16566 -24417
rect 17279 -24397 17313 -24359
rect 17279 -24469 17313 -24431
rect 16396 -24497 16430 -24481
rect 16396 -24569 16430 -24531
rect 14423 -24643 14557 -24627
rect 14423 -24677 14437 -24643
rect 14471 -24677 14509 -24643
rect 14543 -24677 14557 -24643
rect 14423 -24693 14557 -24677
rect 15223 -24647 15493 -24631
rect 15223 -24681 15233 -24647
rect 15267 -24681 15305 -24647
rect 15339 -24681 15377 -24647
rect 15411 -24681 15449 -24647
rect 15483 -24681 15493 -24647
rect 15223 -24699 15493 -24681
rect 16396 -24641 16430 -24603
rect 16396 -24713 16430 -24675
rect 14387 -24773 14421 -24732
rect 13653 -24815 13787 -24799
rect 13653 -24849 13667 -24815
rect 13701 -24849 13739 -24815
rect 13773 -24849 13787 -24815
rect 13653 -24867 13787 -24849
rect 14387 -24845 14421 -24807
rect 13617 -24929 13651 -24913
rect 13617 -25001 13651 -24963
rect 13617 -25051 13651 -25035
rect 13703 -25051 13737 -24913
rect 13789 -24929 13823 -24913
rect 13789 -25001 13823 -24963
rect 13789 -25051 13823 -25035
rect 14387 -24917 14421 -24879
rect 14387 -24989 14421 -24951
rect 14387 -25066 14421 -25023
rect 14473 -25066 14507 -24732
rect 14559 -24773 14593 -24732
rect 14559 -24845 14593 -24807
rect 14559 -24917 14593 -24879
rect 14559 -24989 14593 -24951
rect 14559 -25066 14593 -25023
rect 15169 -24773 15203 -24745
rect 15169 -24845 15203 -24807
rect 15169 -24917 15203 -24879
rect 15169 -24989 15203 -24951
rect 15169 -25051 15203 -25023
rect 15255 -25051 15289 -24745
rect 15341 -24773 15375 -24745
rect 15341 -24845 15375 -24807
rect 15341 -24917 15375 -24879
rect 15341 -24989 15375 -24951
rect 15341 -25051 15375 -25023
rect 15427 -25051 15461 -24745
rect 15513 -24773 15547 -24745
rect 15513 -24845 15547 -24807
rect 15513 -24917 15547 -24879
rect 15513 -24989 15547 -24951
rect 15513 -25051 15547 -25023
rect 16396 -24785 16430 -24747
rect 16396 -24857 16430 -24819
rect 16396 -24929 16430 -24891
rect 16396 -25001 16430 -24963
rect 16396 -25055 16430 -25035
rect 16482 -25051 16516 -24481
rect 16568 -24497 16602 -24481
rect 16568 -24569 16602 -24531
rect 16568 -24641 16602 -24603
rect 16568 -24713 16602 -24675
rect 16568 -24785 16602 -24747
rect 16568 -24857 16602 -24819
rect 16568 -24929 16602 -24891
rect 16568 -25001 16602 -24963
rect 16568 -25051 16602 -25035
rect 17279 -24541 17313 -24503
rect 17279 -24613 17313 -24575
rect 17279 -24685 17313 -24647
rect 17279 -24757 17313 -24719
rect 17279 -24829 17313 -24791
rect 17279 -24901 17313 -24863
rect 17279 -24973 17313 -24935
rect 17279 -25058 17313 -25007
rect 17365 -25058 17399 -24060
rect 17451 -24109 17485 -24060
rect 17451 -24181 17485 -24143
rect 17451 -24253 17485 -24215
rect 17451 -24325 17485 -24287
rect 17451 -24397 17485 -24359
rect 17451 -24469 17485 -24431
rect 17451 -24541 17485 -24503
rect 17451 -24613 17485 -24575
rect 17451 -24685 17485 -24647
rect 17451 -24757 17485 -24719
rect 17451 -24829 17485 -24791
rect 17451 -24901 17485 -24863
rect 17451 -24973 17485 -24935
rect 17451 -25058 17485 -25007
<< obsli1c >>
rect 17377 20625 17411 20659
rect 17449 20625 17483 20659
rect 18089 20625 18123 20659
rect 18161 20625 18195 20659
rect 18233 20625 18267 20659
rect 18305 20625 18339 20659
rect 18917 20625 18951 20659
rect 18989 20625 19023 20659
rect 19061 20625 19095 20659
rect 19133 20625 19167 20659
rect 19205 20625 19239 20659
rect 19277 20625 19311 20659
rect 19349 20625 19383 20659
rect 19421 20625 19455 20659
rect 17327 20513 17361 20547
rect 17327 20441 17361 20475
rect 17327 20369 17361 20403
rect 17327 20297 17361 20331
rect 14889 20193 14923 20227
rect 14961 20193 14995 20227
rect 15447 20193 15481 20227
rect 15519 20193 15553 20227
rect 15591 20193 15625 20227
rect 15663 20193 15697 20227
rect 16118 20193 16152 20227
rect 16190 20193 16224 20227
rect 16262 20193 16296 20227
rect 16334 20193 16368 20227
rect 16406 20193 16440 20227
rect 16478 20193 16512 20227
rect 16550 20193 16584 20227
rect 16622 20193 16656 20227
rect 17327 20225 17361 20259
rect 13865 20109 13899 20143
rect 13937 20109 13971 20143
rect 17327 20153 17361 20187
rect 14839 20081 14873 20115
rect 13815 20009 13849 20043
rect 13987 20009 14021 20043
rect 14839 20009 14873 20043
rect 15011 20081 15045 20115
rect 15011 20009 15045 20043
rect 15383 20081 15417 20115
rect 15383 20009 15417 20043
rect 15555 20081 15589 20115
rect 15555 20009 15589 20043
rect 15727 20081 15761 20115
rect 15727 20009 15761 20043
rect 16026 20081 16060 20115
rect 16026 20009 16060 20043
rect 16198 20081 16232 20115
rect 16198 20009 16232 20043
rect 16370 20081 16404 20115
rect 16370 20009 16404 20043
rect 16542 20081 16576 20115
rect 16542 20009 16576 20043
rect 16714 20081 16748 20115
rect 16714 20009 16748 20043
rect 17327 20081 17361 20115
rect 17327 20009 17361 20043
rect 17499 20513 17533 20547
rect 17499 20441 17533 20475
rect 17499 20369 17533 20403
rect 17499 20297 17533 20331
rect 17499 20225 17533 20259
rect 17499 20153 17533 20187
rect 17499 20081 17533 20115
rect 17499 20009 17533 20043
rect 18025 20513 18059 20547
rect 18025 20441 18059 20475
rect 18025 20369 18059 20403
rect 18025 20297 18059 20331
rect 18025 20225 18059 20259
rect 18025 20153 18059 20187
rect 18025 20081 18059 20115
rect 18025 20009 18059 20043
rect 18197 20513 18231 20547
rect 18197 20441 18231 20475
rect 18197 20369 18231 20403
rect 18197 20297 18231 20331
rect 18197 20225 18231 20259
rect 18197 20153 18231 20187
rect 18197 20081 18231 20115
rect 18197 20009 18231 20043
rect 18369 20513 18403 20547
rect 18369 20441 18403 20475
rect 18369 20369 18403 20403
rect 18369 20297 18403 20331
rect 18369 20225 18403 20259
rect 18369 20153 18403 20187
rect 18369 20081 18403 20115
rect 18369 20009 18403 20043
rect 18825 20513 18859 20547
rect 18825 20441 18859 20475
rect 18825 20369 18859 20403
rect 18825 20297 18859 20331
rect 18825 20225 18859 20259
rect 18825 20153 18859 20187
rect 18825 20081 18859 20115
rect 18825 20009 18859 20043
rect 18997 20513 19031 20547
rect 18997 20441 19031 20475
rect 18997 20369 19031 20403
rect 18997 20297 19031 20331
rect 18997 20225 19031 20259
rect 18997 20153 19031 20187
rect 18997 20081 19031 20115
rect 18997 20009 19031 20043
rect 19169 20513 19203 20547
rect 19169 20441 19203 20475
rect 19169 20369 19203 20403
rect 19169 20297 19203 20331
rect 19169 20225 19203 20259
rect 19169 20153 19203 20187
rect 19169 20081 19203 20115
rect 19169 20009 19203 20043
rect 19341 20513 19375 20547
rect 19341 20441 19375 20475
rect 19341 20369 19375 20403
rect 19341 20297 19375 20331
rect 19341 20225 19375 20259
rect 19341 20153 19375 20187
rect 19341 20081 19375 20115
rect 19341 20009 19375 20043
rect 19513 20513 19547 20547
rect 19513 20441 19547 20475
rect 19513 20369 19547 20403
rect 19513 20297 19547 20331
rect 19513 20225 19547 20259
rect 19513 20153 19547 20187
rect 19513 20081 19547 20115
rect 19513 20009 19547 20043
rect 17329 -24010 17363 -23976
rect 17401 -24010 17435 -23976
rect 17279 -24143 17313 -24109
rect 17279 -24215 17313 -24181
rect 17279 -24287 17313 -24253
rect 17279 -24359 17313 -24325
rect 16446 -24417 16480 -24383
rect 16518 -24417 16552 -24383
rect 17279 -24431 17313 -24397
rect 16396 -24531 16430 -24497
rect 16396 -24603 16430 -24569
rect 14437 -24677 14471 -24643
rect 14509 -24677 14543 -24643
rect 15233 -24681 15267 -24647
rect 15305 -24681 15339 -24647
rect 15377 -24681 15411 -24647
rect 15449 -24681 15483 -24647
rect 16396 -24675 16430 -24641
rect 13667 -24849 13701 -24815
rect 13739 -24849 13773 -24815
rect 14387 -24807 14421 -24773
rect 14387 -24879 14421 -24845
rect 13617 -24963 13651 -24929
rect 13617 -25035 13651 -25001
rect 13789 -24963 13823 -24929
rect 13789 -25035 13823 -25001
rect 14387 -24951 14421 -24917
rect 14387 -25023 14421 -24989
rect 14559 -24807 14593 -24773
rect 14559 -24879 14593 -24845
rect 14559 -24951 14593 -24917
rect 14559 -25023 14593 -24989
rect 15169 -24807 15203 -24773
rect 15169 -24879 15203 -24845
rect 15169 -24951 15203 -24917
rect 15169 -25023 15203 -24989
rect 15341 -24807 15375 -24773
rect 15341 -24879 15375 -24845
rect 15341 -24951 15375 -24917
rect 15341 -25023 15375 -24989
rect 15513 -24807 15547 -24773
rect 15513 -24879 15547 -24845
rect 15513 -24951 15547 -24917
rect 15513 -25023 15547 -24989
rect 16396 -24747 16430 -24713
rect 16396 -24819 16430 -24785
rect 16396 -24891 16430 -24857
rect 16396 -24963 16430 -24929
rect 16396 -25035 16430 -25001
rect 16568 -24531 16602 -24497
rect 16568 -24603 16602 -24569
rect 16568 -24675 16602 -24641
rect 16568 -24747 16602 -24713
rect 16568 -24819 16602 -24785
rect 16568 -24891 16602 -24857
rect 16568 -24963 16602 -24929
rect 16568 -25035 16602 -25001
rect 17279 -24503 17313 -24469
rect 17279 -24575 17313 -24541
rect 17279 -24647 17313 -24613
rect 17279 -24719 17313 -24685
rect 17279 -24791 17313 -24757
rect 17279 -24863 17313 -24829
rect 17279 -24935 17313 -24901
rect 17279 -25007 17313 -24973
rect 17451 -24143 17485 -24109
rect 17451 -24215 17485 -24181
rect 17451 -24287 17485 -24253
rect 17451 -24359 17485 -24325
rect 17451 -24431 17485 -24397
rect 17451 -24503 17485 -24469
rect 17451 -24575 17485 -24541
rect 17451 -24647 17485 -24613
rect 17451 -24719 17485 -24685
rect 17451 -24791 17485 -24757
rect 17451 -24863 17485 -24829
rect 17451 -24935 17485 -24901
rect 17451 -25007 17485 -24973
<< metal1 >>
rect 16968 20659 19467 20671
rect 16968 20625 17377 20659
rect 17411 20625 17449 20659
rect 17483 20625 18089 20659
rect 18123 20625 18161 20659
rect 18195 20625 18233 20659
rect 18267 20625 18305 20659
rect 18339 20625 18917 20659
rect 18951 20625 18989 20659
rect 19023 20625 19061 20659
rect 19095 20625 19133 20659
rect 19167 20625 19205 20659
rect 19239 20625 19277 20659
rect 19311 20625 19349 20659
rect 19383 20625 19421 20659
rect 19455 20625 19467 20659
rect 16968 20613 19467 20625
rect 16968 20239 17042 20613
rect 14436 20227 17042 20239
rect 14436 20193 14889 20227
rect 14923 20193 14961 20227
rect 14995 20193 15447 20227
rect 15481 20193 15519 20227
rect 15553 20193 15591 20227
rect 15625 20193 15663 20227
rect 15697 20193 16118 20227
rect 16152 20193 16190 20227
rect 16224 20193 16262 20227
rect 16296 20193 16334 20227
rect 16368 20193 16406 20227
rect 16440 20193 16478 20227
rect 16512 20193 16550 20227
rect 16584 20193 16622 20227
rect 16656 20193 17042 20227
rect 14436 20181 17042 20193
rect 17321 20547 17367 20563
rect 17321 20513 17327 20547
rect 17361 20513 17367 20547
rect 17321 20475 17367 20513
rect 17321 20441 17327 20475
rect 17361 20441 17367 20475
rect 17321 20403 17367 20441
rect 17321 20369 17327 20403
rect 17361 20369 17367 20403
rect 17321 20331 17367 20369
rect 17321 20297 17327 20331
rect 17361 20297 17367 20331
rect 17321 20259 17367 20297
rect 17321 20225 17327 20259
rect 17361 20225 17367 20259
rect 17321 20187 17367 20225
rect 14436 20157 14510 20181
rect 13652 20143 14510 20157
rect 13652 20109 13865 20143
rect 13899 20109 13937 20143
rect 13971 20109 14510 20143
rect 17321 20153 17327 20187
rect 17361 20153 17367 20187
rect 13652 20097 14510 20109
rect 14833 20115 14879 20131
rect 14833 20081 14839 20115
rect 14873 20081 14879 20115
rect 13809 20043 13855 20062
rect 13809 20009 13815 20043
rect 13849 20009 13855 20043
rect 13809 19913 13855 20009
rect 13981 20043 14027 20062
rect 13981 20009 13987 20043
rect 14021 20009 14027 20043
rect 13981 19913 14027 20009
rect 14833 20043 14879 20081
rect 14833 20009 14839 20043
rect 14873 20009 14879 20043
rect 14833 19913 14879 20009
rect 15005 20115 15051 20131
rect 15005 20081 15011 20115
rect 15045 20081 15051 20115
rect 15005 20043 15051 20081
rect 15005 20009 15011 20043
rect 15045 20009 15051 20043
rect 15005 19913 15051 20009
rect 15377 20115 15423 20131
rect 15377 20081 15383 20115
rect 15417 20081 15423 20115
rect 15377 20043 15423 20081
rect 15377 20009 15383 20043
rect 15417 20009 15423 20043
rect 15377 19913 15423 20009
rect 15549 20115 15595 20131
rect 15549 20081 15555 20115
rect 15589 20081 15595 20115
rect 15549 20043 15595 20081
rect 15549 20009 15555 20043
rect 15589 20009 15595 20043
rect 15549 19913 15595 20009
rect 15721 20115 15767 20131
rect 15721 20081 15727 20115
rect 15761 20081 15767 20115
rect 15721 20043 15767 20081
rect 15721 20009 15727 20043
rect 15761 20009 15767 20043
rect 15721 19913 15767 20009
rect 16020 20115 16066 20131
rect 16020 20081 16026 20115
rect 16060 20081 16066 20115
rect 16020 20043 16066 20081
rect 16020 20009 16026 20043
rect 16060 20009 16066 20043
rect 16020 19913 16066 20009
rect 16192 20115 16238 20131
rect 16192 20081 16198 20115
rect 16232 20081 16238 20115
rect 16192 20043 16238 20081
rect 16192 20009 16198 20043
rect 16232 20009 16238 20043
rect 16192 19913 16238 20009
rect 16364 20115 16410 20131
rect 16364 20081 16370 20115
rect 16404 20081 16410 20115
rect 16364 20043 16410 20081
rect 16364 20009 16370 20043
rect 16404 20009 16410 20043
rect 16364 19913 16410 20009
rect 16536 20115 16582 20131
rect 16536 20081 16542 20115
rect 16576 20081 16582 20115
rect 16536 20043 16582 20081
rect 16536 20009 16542 20043
rect 16576 20009 16582 20043
rect 16536 19913 16582 20009
rect 16708 20115 16754 20131
rect 16708 20081 16714 20115
rect 16748 20081 16754 20115
rect 16708 20043 16754 20081
rect 16708 20009 16714 20043
rect 16748 20009 16754 20043
rect 16708 19913 16754 20009
rect 17321 20115 17367 20153
rect 17321 20081 17327 20115
rect 17361 20081 17367 20115
rect 17321 20043 17367 20081
rect 17321 20009 17327 20043
rect 17361 20009 17367 20043
rect 17321 19913 17367 20009
rect 17493 20547 17539 20563
rect 17493 20513 17499 20547
rect 17533 20513 17539 20547
rect 17493 20475 17539 20513
rect 17493 20441 17499 20475
rect 17533 20441 17539 20475
rect 17493 20403 17539 20441
rect 17493 20369 17499 20403
rect 17533 20369 17539 20403
rect 17493 20331 17539 20369
rect 17493 20297 17499 20331
rect 17533 20297 17539 20331
rect 17493 20259 17539 20297
rect 17493 20225 17499 20259
rect 17533 20225 17539 20259
rect 17493 20187 17539 20225
rect 17493 20153 17499 20187
rect 17533 20153 17539 20187
rect 17493 20115 17539 20153
rect 17493 20081 17499 20115
rect 17533 20081 17539 20115
rect 17493 20043 17539 20081
rect 17493 20009 17499 20043
rect 17533 20009 17539 20043
rect 17493 19913 17539 20009
rect 18019 20547 18065 20563
rect 18019 20513 18025 20547
rect 18059 20513 18065 20547
rect 18019 20475 18065 20513
rect 18019 20441 18025 20475
rect 18059 20441 18065 20475
rect 18019 20403 18065 20441
rect 18019 20369 18025 20403
rect 18059 20369 18065 20403
rect 18019 20331 18065 20369
rect 18019 20297 18025 20331
rect 18059 20297 18065 20331
rect 18019 20259 18065 20297
rect 18019 20225 18025 20259
rect 18059 20225 18065 20259
rect 18019 20187 18065 20225
rect 18019 20153 18025 20187
rect 18059 20153 18065 20187
rect 18019 20115 18065 20153
rect 18019 20081 18025 20115
rect 18059 20081 18065 20115
rect 18019 20043 18065 20081
rect 18019 20009 18025 20043
rect 18059 20009 18065 20043
rect 18019 19913 18065 20009
rect 18191 20547 18237 20563
rect 18191 20513 18197 20547
rect 18231 20513 18237 20547
rect 18191 20475 18237 20513
rect 18191 20441 18197 20475
rect 18231 20441 18237 20475
rect 18191 20403 18237 20441
rect 18191 20369 18197 20403
rect 18231 20369 18237 20403
rect 18191 20331 18237 20369
rect 18191 20297 18197 20331
rect 18231 20297 18237 20331
rect 18191 20259 18237 20297
rect 18191 20225 18197 20259
rect 18231 20225 18237 20259
rect 18191 20187 18237 20225
rect 18191 20153 18197 20187
rect 18231 20153 18237 20187
rect 18191 20115 18237 20153
rect 18191 20081 18197 20115
rect 18231 20081 18237 20115
rect 18191 20043 18237 20081
rect 18191 20009 18197 20043
rect 18231 20009 18237 20043
rect 18191 19913 18237 20009
rect 18363 20547 18409 20563
rect 18363 20513 18369 20547
rect 18403 20513 18409 20547
rect 18363 20475 18409 20513
rect 18363 20441 18369 20475
rect 18403 20441 18409 20475
rect 18363 20403 18409 20441
rect 18363 20369 18369 20403
rect 18403 20369 18409 20403
rect 18363 20331 18409 20369
rect 18363 20297 18369 20331
rect 18403 20297 18409 20331
rect 18363 20259 18409 20297
rect 18363 20225 18369 20259
rect 18403 20225 18409 20259
rect 18363 20187 18409 20225
rect 18363 20153 18369 20187
rect 18403 20153 18409 20187
rect 18363 20115 18409 20153
rect 18363 20081 18369 20115
rect 18403 20081 18409 20115
rect 18363 20043 18409 20081
rect 18363 20009 18369 20043
rect 18403 20009 18409 20043
rect 18363 19913 18409 20009
rect 18819 20547 18865 20563
rect 18819 20513 18825 20547
rect 18859 20513 18865 20547
rect 18819 20475 18865 20513
rect 18819 20441 18825 20475
rect 18859 20441 18865 20475
rect 18819 20403 18865 20441
rect 18819 20369 18825 20403
rect 18859 20369 18865 20403
rect 18819 20331 18865 20369
rect 18819 20297 18825 20331
rect 18859 20297 18865 20331
rect 18819 20259 18865 20297
rect 18819 20225 18825 20259
rect 18859 20225 18865 20259
rect 18819 20187 18865 20225
rect 18819 20153 18825 20187
rect 18859 20153 18865 20187
rect 18819 20115 18865 20153
rect 18819 20081 18825 20115
rect 18859 20081 18865 20115
rect 18819 20043 18865 20081
rect 18819 20009 18825 20043
rect 18859 20009 18865 20043
rect 18819 19913 18865 20009
rect 18991 20547 19037 20563
rect 18991 20513 18997 20547
rect 19031 20513 19037 20547
rect 18991 20475 19037 20513
rect 18991 20441 18997 20475
rect 19031 20441 19037 20475
rect 18991 20403 19037 20441
rect 18991 20369 18997 20403
rect 19031 20369 19037 20403
rect 18991 20331 19037 20369
rect 18991 20297 18997 20331
rect 19031 20297 19037 20331
rect 18991 20259 19037 20297
rect 18991 20225 18997 20259
rect 19031 20225 19037 20259
rect 18991 20187 19037 20225
rect 18991 20153 18997 20187
rect 19031 20153 19037 20187
rect 18991 20115 19037 20153
rect 18991 20081 18997 20115
rect 19031 20081 19037 20115
rect 18991 20043 19037 20081
rect 18991 20009 18997 20043
rect 19031 20009 19037 20043
rect 18991 19913 19037 20009
rect 19163 20547 19209 20563
rect 19163 20513 19169 20547
rect 19203 20513 19209 20547
rect 19163 20475 19209 20513
rect 19163 20441 19169 20475
rect 19203 20441 19209 20475
rect 19163 20403 19209 20441
rect 19163 20369 19169 20403
rect 19203 20369 19209 20403
rect 19163 20331 19209 20369
rect 19163 20297 19169 20331
rect 19203 20297 19209 20331
rect 19163 20259 19209 20297
rect 19163 20225 19169 20259
rect 19203 20225 19209 20259
rect 19163 20187 19209 20225
rect 19163 20153 19169 20187
rect 19203 20153 19209 20187
rect 19163 20115 19209 20153
rect 19163 20081 19169 20115
rect 19203 20081 19209 20115
rect 19163 20043 19209 20081
rect 19163 20009 19169 20043
rect 19203 20009 19209 20043
rect 19163 19913 19209 20009
rect 19335 20547 19381 20563
rect 19335 20513 19341 20547
rect 19375 20513 19381 20547
rect 19335 20475 19381 20513
rect 19335 20441 19341 20475
rect 19375 20441 19381 20475
rect 19335 20403 19381 20441
rect 19335 20369 19341 20403
rect 19375 20369 19381 20403
rect 19335 20331 19381 20369
rect 19335 20297 19341 20331
rect 19375 20297 19381 20331
rect 19335 20259 19381 20297
rect 19335 20225 19341 20259
rect 19375 20225 19381 20259
rect 19335 20187 19381 20225
rect 19335 20153 19341 20187
rect 19375 20153 19381 20187
rect 19335 20115 19381 20153
rect 19335 20081 19341 20115
rect 19375 20081 19381 20115
rect 19335 20043 19381 20081
rect 19335 20009 19341 20043
rect 19375 20009 19381 20043
rect 19335 19913 19381 20009
rect 19507 20547 19553 20563
rect 19507 20513 19513 20547
rect 19547 20513 19553 20547
rect 19507 20475 19553 20513
rect 19507 20441 19513 20475
rect 19547 20441 19553 20475
rect 19507 20403 19553 20441
rect 19507 20369 19513 20403
rect 19547 20369 19553 20403
rect 19507 20331 19553 20369
rect 19507 20297 19513 20331
rect 19547 20297 19553 20331
rect 19507 20259 19553 20297
rect 19507 20225 19513 20259
rect 19547 20225 19553 20259
rect 19507 20187 19553 20225
rect 19507 20153 19513 20187
rect 19547 20153 19553 20187
rect 19507 20115 19553 20153
rect 19507 20081 19513 20115
rect 19547 20081 19553 20115
rect 19507 20043 19553 20081
rect 19507 20009 19513 20043
rect 19547 20009 19553 20043
rect 19507 19913 19553 20009
rect 13652 19853 19553 19913
rect 16941 -23976 17447 -23964
rect 16941 -24010 17329 -23976
rect 17363 -24010 17401 -23976
rect 17435 -24010 17447 -23976
rect 16941 -24022 17447 -24010
rect 16941 -24371 17010 -24022
rect 15875 -24383 17010 -24371
rect 15875 -24417 16446 -24383
rect 16480 -24417 16518 -24383
rect 16552 -24417 17010 -24383
rect 15875 -24429 17010 -24417
rect 17273 -24109 17319 -24060
rect 17273 -24143 17279 -24109
rect 17313 -24143 17319 -24109
rect 17273 -24181 17319 -24143
rect 17273 -24215 17279 -24181
rect 17313 -24215 17319 -24181
rect 17273 -24253 17319 -24215
rect 17273 -24287 17279 -24253
rect 17313 -24287 17319 -24253
rect 17273 -24325 17319 -24287
rect 17273 -24359 17279 -24325
rect 17313 -24359 17319 -24325
rect 17273 -24397 17319 -24359
rect 15875 -24631 15944 -24429
rect 17273 -24431 17279 -24397
rect 17313 -24431 17319 -24397
rect 17273 -24469 17319 -24431
rect 14089 -24643 15944 -24631
rect 14089 -24677 14437 -24643
rect 14471 -24677 14509 -24643
rect 14543 -24647 15944 -24643
rect 14543 -24677 15233 -24647
rect 14089 -24681 15233 -24677
rect 15267 -24681 15305 -24647
rect 15339 -24681 15377 -24647
rect 15411 -24681 15449 -24647
rect 15483 -24681 15944 -24647
rect 14089 -24689 15944 -24681
rect 16390 -24497 16436 -24481
rect 16390 -24531 16396 -24497
rect 16430 -24531 16436 -24497
rect 16390 -24569 16436 -24531
rect 16390 -24603 16396 -24569
rect 16430 -24603 16436 -24569
rect 16390 -24641 16436 -24603
rect 16390 -24675 16396 -24641
rect 16430 -24675 16436 -24641
rect 14089 -24803 14158 -24689
rect 15221 -24693 15495 -24689
rect 16390 -24713 16436 -24675
rect 13326 -24815 14158 -24803
rect 13326 -24849 13667 -24815
rect 13701 -24849 13739 -24815
rect 13773 -24849 14158 -24815
rect 13326 -24861 14158 -24849
rect 14381 -24773 14427 -24732
rect 14381 -24807 14387 -24773
rect 14421 -24807 14427 -24773
rect 14381 -24845 14427 -24807
rect 14381 -24879 14387 -24845
rect 14421 -24879 14427 -24845
rect 13611 -24929 13657 -24913
rect 13611 -24963 13617 -24929
rect 13651 -24963 13657 -24929
rect 13611 -25001 13657 -24963
rect 13611 -25035 13617 -25001
rect 13651 -25035 13657 -25001
rect 13611 -25131 13657 -25035
rect 13783 -24929 13829 -24913
rect 13783 -24963 13789 -24929
rect 13823 -24963 13829 -24929
rect 13783 -25001 13829 -24963
rect 13783 -25035 13789 -25001
rect 13823 -25035 13829 -25001
rect 13783 -25131 13829 -25035
rect 14381 -24917 14427 -24879
rect 14381 -24951 14387 -24917
rect 14421 -24951 14427 -24917
rect 14381 -24989 14427 -24951
rect 14381 -25023 14387 -24989
rect 14421 -25023 14427 -24989
rect 14381 -25131 14427 -25023
rect 14553 -24773 14599 -24732
rect 14553 -24807 14559 -24773
rect 14593 -24807 14599 -24773
rect 14553 -24845 14599 -24807
rect 14553 -24879 14559 -24845
rect 14593 -24879 14599 -24845
rect 14553 -24917 14599 -24879
rect 14553 -24951 14559 -24917
rect 14593 -24951 14599 -24917
rect 14553 -24989 14599 -24951
rect 14553 -25023 14559 -24989
rect 14593 -25023 14599 -24989
rect 14553 -25131 14599 -25023
rect 15163 -24773 15209 -24745
rect 15163 -24807 15169 -24773
rect 15203 -24807 15209 -24773
rect 15163 -24845 15209 -24807
rect 15163 -24879 15169 -24845
rect 15203 -24879 15209 -24845
rect 15163 -24917 15209 -24879
rect 15163 -24951 15169 -24917
rect 15203 -24951 15209 -24917
rect 15163 -24989 15209 -24951
rect 15163 -25023 15169 -24989
rect 15203 -25023 15209 -24989
rect 15163 -25131 15209 -25023
rect 15335 -24773 15381 -24745
rect 15335 -24807 15341 -24773
rect 15375 -24807 15381 -24773
rect 15335 -24845 15381 -24807
rect 15335 -24879 15341 -24845
rect 15375 -24879 15381 -24845
rect 15335 -24917 15381 -24879
rect 15335 -24951 15341 -24917
rect 15375 -24951 15381 -24917
rect 15335 -24989 15381 -24951
rect 15335 -25023 15341 -24989
rect 15375 -25023 15381 -24989
rect 15335 -25131 15381 -25023
rect 15507 -24773 15553 -24745
rect 15507 -24807 15513 -24773
rect 15547 -24807 15553 -24773
rect 15507 -24845 15553 -24807
rect 15507 -24879 15513 -24845
rect 15547 -24879 15553 -24845
rect 15507 -24917 15553 -24879
rect 15507 -24951 15513 -24917
rect 15547 -24951 15553 -24917
rect 15507 -24989 15553 -24951
rect 15507 -25023 15513 -24989
rect 15547 -25023 15553 -24989
rect 15507 -25131 15553 -25023
rect 16390 -24747 16396 -24713
rect 16430 -24747 16436 -24713
rect 16390 -24785 16436 -24747
rect 16390 -24819 16396 -24785
rect 16430 -24819 16436 -24785
rect 16390 -24857 16436 -24819
rect 16390 -24891 16396 -24857
rect 16430 -24891 16436 -24857
rect 16390 -24929 16436 -24891
rect 16390 -24963 16396 -24929
rect 16430 -24963 16436 -24929
rect 16390 -25001 16436 -24963
rect 16390 -25035 16396 -25001
rect 16430 -25035 16436 -25001
rect 16390 -25131 16436 -25035
rect 16562 -24497 16608 -24481
rect 16562 -24531 16568 -24497
rect 16602 -24531 16608 -24497
rect 16562 -24569 16608 -24531
rect 16562 -24603 16568 -24569
rect 16602 -24603 16608 -24569
rect 16562 -24641 16608 -24603
rect 16562 -24675 16568 -24641
rect 16602 -24675 16608 -24641
rect 16562 -24713 16608 -24675
rect 16562 -24747 16568 -24713
rect 16602 -24747 16608 -24713
rect 16562 -24785 16608 -24747
rect 16562 -24819 16568 -24785
rect 16602 -24819 16608 -24785
rect 16562 -24857 16608 -24819
rect 16562 -24891 16568 -24857
rect 16602 -24891 16608 -24857
rect 16562 -24929 16608 -24891
rect 16562 -24963 16568 -24929
rect 16602 -24963 16608 -24929
rect 16562 -25001 16608 -24963
rect 16562 -25035 16568 -25001
rect 16602 -25035 16608 -25001
rect 16562 -25131 16608 -25035
rect 17273 -24503 17279 -24469
rect 17313 -24503 17319 -24469
rect 17273 -24541 17319 -24503
rect 17273 -24575 17279 -24541
rect 17313 -24575 17319 -24541
rect 17273 -24613 17319 -24575
rect 17273 -24647 17279 -24613
rect 17313 -24647 17319 -24613
rect 17273 -24685 17319 -24647
rect 17273 -24719 17279 -24685
rect 17313 -24719 17319 -24685
rect 17273 -24757 17319 -24719
rect 17273 -24791 17279 -24757
rect 17313 -24791 17319 -24757
rect 17273 -24829 17319 -24791
rect 17273 -24863 17279 -24829
rect 17313 -24863 17319 -24829
rect 17273 -24901 17319 -24863
rect 17273 -24935 17279 -24901
rect 17313 -24935 17319 -24901
rect 17273 -24973 17319 -24935
rect 17273 -25007 17279 -24973
rect 17313 -25007 17319 -24973
rect 17273 -25131 17319 -25007
rect 17445 -24109 17491 -24060
rect 17445 -24143 17451 -24109
rect 17485 -24143 17491 -24109
rect 17445 -24181 17491 -24143
rect 17445 -24215 17451 -24181
rect 17485 -24215 17491 -24181
rect 17445 -24253 17491 -24215
rect 17445 -24287 17451 -24253
rect 17485 -24287 17491 -24253
rect 17445 -24325 17491 -24287
rect 17445 -24359 17451 -24325
rect 17485 -24359 17491 -24325
rect 17445 -24397 17491 -24359
rect 17445 -24431 17451 -24397
rect 17485 -24431 17491 -24397
rect 17445 -24469 17491 -24431
rect 17445 -24503 17451 -24469
rect 17485 -24503 17491 -24469
rect 17445 -24541 17491 -24503
rect 17445 -24575 17451 -24541
rect 17485 -24575 17491 -24541
rect 17445 -24613 17491 -24575
rect 17445 -24647 17451 -24613
rect 17485 -24647 17491 -24613
rect 17445 -24685 17491 -24647
rect 17445 -24719 17451 -24685
rect 17485 -24719 17491 -24685
rect 17445 -24757 17491 -24719
rect 17445 -24791 17451 -24757
rect 17485 -24791 17491 -24757
rect 17445 -24829 17491 -24791
rect 17445 -24863 17451 -24829
rect 17485 -24863 17491 -24829
rect 17445 -24901 17491 -24863
rect 17445 -24935 17451 -24901
rect 17485 -24935 17491 -24901
rect 17445 -24973 17491 -24935
rect 17445 -25007 17451 -24973
rect 17485 -25007 17491 -24973
rect 17445 -25131 17491 -25007
rect 13326 -25191 17491 -25131
<< obsm1 >>
rect 13892 19993 13944 20062
rect 14916 19993 14968 20131
rect 15460 19993 15512 20131
rect 15632 19993 15684 20131
rect 16103 19993 16155 20131
rect 16275 19993 16327 20131
rect 16447 19993 16499 20131
rect 16619 19993 16671 20131
rect 17404 19993 17456 20563
rect 18102 19993 18154 20563
rect 18274 19993 18326 20563
rect 18902 19993 18954 20563
rect 19074 19993 19126 20563
rect 19246 19993 19298 20563
rect 19418 19993 19470 20563
rect 13694 -25051 13746 -24913
rect 14464 -25066 14516 -24732
rect 15246 -25051 15298 -24745
rect 15418 -25051 15470 -24745
rect 16473 -25051 16525 -24481
rect 17356 -25058 17408 -24060
<< obsm2 >>
rect 17166 20430 17858 20575
rect 18095 20415 18161 20569
rect 18267 20415 18333 20569
rect 18895 20415 18961 20569
rect 19067 20415 19133 20569
rect 19239 20415 19305 20569
rect 19411 20415 19477 20569
rect 14916 20062 14968 20126
rect 13652 19993 15260 20062
rect 15453 19983 15519 20137
rect 15625 19983 15691 20137
rect 16096 19983 16162 20137
rect 16268 19983 16334 20137
rect 16440 19983 16506 20137
rect 16612 19983 16678 20137
rect 17061 -24190 17408 -24062
rect 17061 -24486 17170 -24190
rect 16068 -24614 17170 -24486
rect 14225 -24861 15017 -24733
rect 14225 -24918 14298 -24861
rect 15239 -24891 15305 -24737
rect 15411 -24891 15477 -24737
rect 16068 -24862 16177 -24614
rect 13327 -25046 14298 -24918
<< metal3 >>
rect 17166 20137 17244 20575
rect 17756 20415 19477 20575
rect 15179 19993 17244 20137
rect 15453 19983 15519 19993
rect 15625 19983 15691 19993
rect 16096 19983 16162 19993
rect 16268 19983 16334 19993
rect 16440 19983 16506 19993
rect 16612 19983 16678 19993
rect 14892 -24862 16177 -24733
rect 15239 -24891 15305 -24862
rect 15411 -24891 15477 -24862
<< labels >>
rlabel locali s 1835 -41064 2397 -40469 8 B_P
port 1 nsew
rlabel metal3 s 15411 -24891 15477 -24862 8 D_P
port 2 nsew
rlabel metal3 s 15239 -24891 15305 -24862 8 D_P
port 2 nsew
rlabel metal3 s 14892 -24862 16177 -24733 8 D_P
port 2 nsew
rlabel metal1 s 16968 20613 19467 20671 6 G
port 3 nsew
rlabel metal1 s 16968 20239 17042 20613 6 G
port 3 nsew
rlabel metal1 s 14436 20181 17042 20239 6 G
port 3 nsew
rlabel metal1 s 14436 20157 14510 20181 6 G
port 3 nsew
rlabel metal1 s 13652 20097 14510 20157 6 G
port 3 nsew
rlabel metal1 s 16941 -24022 17447 -23964 8 G_P
port 4 nsew
rlabel metal1 s 16941 -24371 17010 -24022 8 G_P
port 4 nsew
rlabel metal1 s 15875 -24429 17010 -24371 8 G_P
port 4 nsew
rlabel metal1 s 15875 -24631 15944 -24429 8 G_P
port 4 nsew
rlabel metal1 s 15221 -24693 15495 -24689 8 G_P
port 4 nsew
rlabel metal1 s 14089 -24689 15944 -24631 8 G_P
port 4 nsew
rlabel metal1 s 14089 -24803 14158 -24689 8 G_P
port 4 nsew
rlabel metal1 s 13326 -24861 14158 -24803 8 G_P
port 4 nsew
rlabel locali s 1835 1730 2397 2325 6 NWELL
port 5 nsew
rlabel metal1 s 19507 19913 19553 20563 6 S
port 6 nsew
rlabel metal1 s 19335 19913 19381 20563 6 S
port 6 nsew
rlabel metal1 s 19163 19913 19209 20563 6 S
port 6 nsew
rlabel metal1 s 18991 19913 19037 20563 6 S
port 6 nsew
rlabel metal1 s 18819 19913 18865 20563 6 S
port 6 nsew
rlabel metal1 s 18363 19913 18409 20563 6 S
port 6 nsew
rlabel metal1 s 18191 19913 18237 20563 6 S
port 6 nsew
rlabel metal1 s 18019 19913 18065 20563 6 S
port 6 nsew
rlabel metal1 s 17493 19913 17539 20563 6 S
port 6 nsew
rlabel metal1 s 17321 19913 17367 20563 6 S
port 6 nsew
rlabel metal1 s 16708 19913 16754 20131 6 S
port 6 nsew
rlabel metal1 s 16536 19913 16582 20131 6 S
port 6 nsew
rlabel metal1 s 16364 19913 16410 20131 6 S
port 6 nsew
rlabel metal1 s 16192 19913 16238 20131 6 S
port 6 nsew
rlabel metal1 s 16020 19913 16066 20131 6 S
port 6 nsew
rlabel metal1 s 15721 19913 15767 20131 6 S
port 6 nsew
rlabel metal1 s 15549 19913 15595 20131 6 S
port 6 nsew
rlabel metal1 s 15377 19913 15423 20131 6 S
port 6 nsew
rlabel metal1 s 15005 19913 15051 20131 6 S
port 6 nsew
rlabel metal1 s 14833 19913 14879 20131 6 S
port 6 nsew
rlabel metal1 s 13981 19913 14027 20062 6 S
port 6 nsew
rlabel metal1 s 13809 19913 13855 20062 6 S
port 6 nsew
rlabel metal1 s 13652 19853 19553 19913 6 S
port 6 nsew
rlabel metal1 s 17445 -25131 17491 -24060 8 S_P
port 7 nsew
rlabel metal1 s 17273 -25131 17319 -24060 8 S_P
port 7 nsew
rlabel metal1 s 16562 -25131 16608 -24481 8 S_P
port 7 nsew
rlabel metal1 s 16390 -25131 16436 -24481 8 S_P
port 7 nsew
rlabel metal1 s 15507 -25131 15553 -24745 8 S_P
port 7 nsew
rlabel metal1 s 15335 -25131 15381 -24745 8 S_P
port 7 nsew
rlabel metal1 s 15163 -25131 15209 -24745 8 S_P
port 7 nsew
rlabel metal1 s 14553 -25131 14599 -24732 8 S_P
port 7 nsew
rlabel metal1 s 14381 -25131 14427 -24732 8 S_P
port 7 nsew
rlabel metal1 s 13783 -25131 13829 -24913 8 S_P
port 7 nsew
rlabel metal1 s 13611 -25131 13657 -24913 8 S_P
port 7 nsew
rlabel metal1 s 13326 -25191 17491 -25131 8 S_P
port 7 nsew
rlabel locali s 12028 18138 12590 18733 6 VGND
port 8 nsew ground default
rlabel metal3 s 17756 20415 19477 20575 6 VPWR
port 9 nsew power default
rlabel metal3 s 17166 20137 17244 20575 6 VPWR
port 9 nsew power default
rlabel metal3 s 16612 19983 16678 19993 6 VPWR
port 9 nsew power default
rlabel metal3 s 16440 19983 16506 19993 6 VPWR
port 9 nsew power default
rlabel metal3 s 16268 19983 16334 19993 6 VPWR
port 9 nsew power default
rlabel metal3 s 16096 19983 16162 19993 6 VPWR
port 9 nsew power default
rlabel metal3 s 15625 19983 15691 19993 6 VPWR
port 9 nsew power default
rlabel metal3 s 15453 19983 15519 19993 6 VPWR
port 9 nsew power default
rlabel metal3 s 15179 19993 17244 20137 6 VPWR
port 9 nsew power default
<< properties >>
string FIXED_BBOX 0 -42794 311106 39640
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10553276
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10548138
<< end >>
