magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< poly >>
rect -160 10457 0 10473
rect -160 10423 -131 10457
rect -97 10423 -63 10457
rect -29 10423 0 10457
rect -160 10089 -131 10123
rect -97 10089 -63 10123
rect -29 10089 0 10123
rect -160 10073 0 10089
rect 517 10437 677 10453
rect 517 10403 546 10437
rect 580 10403 614 10437
rect 648 10403 677 10437
rect 517 10069 546 10103
rect 580 10069 614 10103
rect 648 10069 677 10103
rect 517 10053 677 10069
rect -160 9872 0 9888
rect -160 9838 -131 9872
rect -97 9838 -63 9872
rect -29 9838 0 9872
rect -160 9504 -131 9538
rect -97 9504 -63 9538
rect -29 9504 0 9538
rect -160 9488 0 9504
rect 517 9852 677 9868
rect 517 9818 546 9852
rect 580 9818 614 9852
rect 648 9818 677 9852
rect 517 9484 546 9518
rect 580 9484 614 9518
rect 648 9484 677 9518
rect 517 9468 677 9484
<< polycont >>
rect -131 10423 -97 10457
rect -63 10423 -29 10457
rect -131 10089 -97 10123
rect -63 10089 -29 10123
rect 546 10403 580 10437
rect 614 10403 648 10437
rect 546 10069 580 10103
rect 614 10069 648 10103
rect -131 9838 -97 9872
rect -63 9838 -29 9872
rect -131 9504 -97 9538
rect -63 9504 -29 9538
rect 546 9818 580 9852
rect 614 9818 648 9852
rect 546 9484 580 9518
rect 614 9484 648 9518
<< npolyres >>
rect -160 10123 0 10423
rect 517 10103 677 10403
rect -160 9538 0 9838
rect 517 9518 677 9818
<< locali >>
rect -147 10430 -133 10536
rect -27 10430 -13 10536
rect -147 10423 -131 10430
rect -97 10423 -63 10430
rect -29 10423 -13 10430
rect 530 10431 544 10537
rect 650 10431 664 10537
rect 530 10403 546 10431
rect 580 10403 614 10431
rect 648 10403 664 10431
rect -147 10102 -131 10123
rect -147 10068 -133 10102
rect -97 10089 -63 10123
rect -29 10102 -13 10123
rect -99 10068 -61 10089
rect -27 10068 -13 10102
rect -147 9974 -13 10068
rect -147 9868 -133 9974
rect -27 9868 -13 9974
rect -147 9838 -131 9868
rect -97 9838 -63 9868
rect -29 9838 -13 9868
rect 530 10069 544 10103
rect 580 10069 614 10103
rect 650 10069 664 10103
rect 530 9985 664 10069
rect 530 9879 544 9985
rect 650 9879 664 9985
rect 530 9852 664 9879
rect 530 9818 546 9852
rect 580 9818 614 9852
rect 648 9818 664 9852
rect -147 9504 -133 9538
rect -97 9504 -63 9538
rect -27 9504 -13 9538
rect 530 9484 544 9518
rect 580 9484 614 9518
rect 650 9484 664 9518
rect -99 9396 -61 9430
rect 578 8772 616 8806
rect -101 8162 -63 8196
rect -101 8054 -63 8088
rect -101 6820 -63 6854
rect 98 6152 410 6158
rect 98 6046 110 6152
rect 216 6046 410 6152
<< viali >>
rect -133 10457 -27 10536
rect -133 10430 -131 10457
rect -131 10430 -97 10457
rect -97 10430 -63 10457
rect -63 10430 -29 10457
rect -29 10430 -27 10457
rect 544 10437 650 10537
rect 544 10431 546 10437
rect 546 10431 580 10437
rect 580 10431 614 10437
rect 614 10431 648 10437
rect 648 10431 650 10437
rect -133 10089 -131 10102
rect -131 10089 -99 10102
rect -61 10089 -29 10102
rect -29 10089 -27 10102
rect -133 10068 -99 10089
rect -61 10068 -27 10089
rect -133 9872 -27 9974
rect -133 9868 -131 9872
rect -131 9868 -97 9872
rect -97 9868 -63 9872
rect -63 9868 -29 9872
rect -29 9868 -27 9872
rect 544 10069 546 10103
rect 546 10069 578 10103
rect 616 10069 648 10103
rect 648 10069 650 10103
rect 544 9879 650 9985
rect -133 9504 -131 9538
rect -131 9504 -99 9538
rect -61 9504 -29 9538
rect -29 9504 -27 9538
rect 544 9484 546 9518
rect 546 9484 578 9518
rect 616 9484 648 9518
rect 648 9484 650 9518
rect -133 9396 -99 9430
rect -61 9396 -27 9430
rect 544 8772 578 8806
rect 616 8772 650 8806
rect -135 8162 -101 8196
rect -63 8162 -29 8196
rect -135 8054 -101 8088
rect -63 8054 -29 8088
rect -135 6820 -101 6854
rect -63 6820 -29 6854
rect 110 6046 216 6152
<< metal1 >>
rect -147 10537 664 10611
rect -147 10536 544 10537
rect -147 10430 -133 10536
rect -27 10483 544 10536
rect -27 10431 -9 10483
tri -9 10431 43 10483 nw
tri 504 10455 532 10483 ne
rect 532 10431 544 10483
rect 650 10431 664 10537
rect -27 10430 -15 10431
rect -147 10417 -15 10430
tri -15 10425 -9 10431 nw
rect -146 10415 -16 10416
rect -147 10115 -15 10415
rect -146 10114 -16 10115
rect -147 10102 -15 10113
rect -147 10068 -133 10102
rect -99 10068 -61 10102
rect -27 10068 -15 10102
rect -147 9974 -15 10068
rect -147 9868 -133 9974
rect -27 9868 -15 9974
rect -147 9857 -15 9868
rect -146 9855 -16 9856
rect -147 9555 -15 9855
rect -146 9554 -16 9555
rect -147 9538 -15 9553
rect -147 9504 -133 9538
rect -99 9504 -61 9538
rect -27 9504 -15 9538
rect -147 9430 -15 9504
rect 532 10417 664 10431
rect 533 10415 663 10416
rect 532 10115 664 10415
rect 533 10114 663 10115
rect 532 10103 664 10113
rect 532 10069 544 10103
rect 578 10069 616 10103
rect 650 10069 664 10103
rect 532 9985 664 10069
rect 532 9879 544 9985
rect 650 9879 664 9985
rect 532 9836 664 9879
rect 533 9834 663 9835
rect 532 9534 664 9834
rect 533 9533 663 9534
rect 532 9518 664 9532
rect 532 9484 544 9518
rect 578 9484 616 9518
rect 650 9484 664 9518
rect 532 9478 664 9484
rect -147 9396 -133 9430
rect -99 9396 -61 9430
rect -27 9396 -15 9430
rect -147 9079 -15 9396
rect -146 9077 -16 9078
rect -147 8777 -15 9077
rect -146 8776 -16 8777
rect -147 8196 -15 8775
rect -147 8162 -135 8196
rect -101 8162 -63 8196
rect -29 8162 -15 8196
rect -147 8088 -15 8162
rect -147 8054 -135 8088
rect -101 8054 -63 8088
rect -29 8054 -15 8088
rect -147 7737 -15 8054
rect -146 7735 -16 7736
rect 532 8806 662 8812
rect 532 8772 544 8806
rect 578 8772 616 8806
rect 650 8772 662 8806
rect -146 7434 -16 7435
rect -147 6860 -15 7433
tri -15 6860 10 6885 sw
tri 507 6860 532 6885 se
rect 532 6860 662 8772
rect -147 6854 662 6860
rect -147 6820 -135 6854
rect -101 6820 -63 6854
rect -29 6820 662 6854
rect -147 6779 662 6820
rect 98 6152 228 6158
rect 98 6046 110 6152
rect 216 6046 228 6152
rect 98 6040 228 6046
<< rmetal1 >>
rect -147 10416 -15 10417
rect -147 10415 -146 10416
rect -16 10415 -15 10416
rect -147 10114 -146 10115
rect -16 10114 -15 10115
rect -147 10113 -15 10114
rect -147 9856 -15 9857
rect -147 9855 -146 9856
rect -16 9855 -15 9856
rect -147 9554 -146 9555
rect -16 9554 -15 9555
rect -147 9553 -15 9554
rect 532 10416 664 10417
rect 532 10415 533 10416
rect 663 10415 664 10416
rect 532 10114 533 10115
rect 663 10114 664 10115
rect 532 10113 664 10114
rect 532 9835 664 9836
rect 532 9834 533 9835
rect 663 9834 664 9835
rect 532 9533 533 9534
rect 663 9533 664 9534
rect 532 9532 664 9533
rect -147 9078 -15 9079
rect -147 9077 -146 9078
rect -16 9077 -15 9078
rect -147 8776 -146 8777
rect -16 8776 -15 8777
rect -147 8775 -15 8776
rect -147 7736 -15 7737
rect -147 7735 -146 7736
rect -16 7735 -15 7736
rect -147 7434 -146 7435
rect -16 7434 -15 7435
rect -147 7433 -15 7434
use sky130_fd_io__com_res_weak_bentbigres  sky130_fd_io__com_res_weak_bentbigres_0
timestamp 1679235063
transform -1 0 421 0 1 0
box -258 1014 579 9446
use sky130_fd_io__tk_em1o_cdns_5595914180860  sky130_fd_io__tk_em1o_cdns_5595914180860_0
timestamp 1679235063
transform 0 -1 -15 1 0 7381
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_0
timestamp 1679235063
transform 0 -1 -15 1 0 8723
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_1
timestamp 1679235063
transform 0 1 532 -1 0 9888
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_2
timestamp 1679235063
transform 0 1 532 -1 0 10469
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_3
timestamp 1679235063
transform 0 -1 -15 1 0 10061
box 0 0 1 1
use sky130_fd_io__tk_em1s_cdns_5595914180859  sky130_fd_io__tk_em1s_cdns_5595914180859_4
timestamp 1679235063
transform 0 -1 -15 1 0 9501
box 0 0 1 1
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_0
timestamp 1679235063
transform 0 1 517 -1 0 9818
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_1
timestamp 1679235063
transform 0 1 517 -1 0 10403
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_2
timestamp 1679235063
transform 0 -1 0 1 0 10123
box 15 13 285 14
use sky130_fd_pr__res_generic_po__example_5595914180864  sky130_fd_pr__res_generic_po__example_5595914180864_3
timestamp 1679235063
transform 0 -1 0 1 0 9538
box 15 13 285 14
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1679235063
transform 1 0 544 0 1 8772
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_1
timestamp 1679235063
transform 1 0 -135 0 1 6820
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_2
timestamp 1679235063
transform 1 0 -135 0 1 8162
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_3
timestamp 1679235063
transform -1 0 -27 0 1 9396
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_4
timestamp 1679235063
transform 1 0 -135 0 1 8054
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_5
timestamp 1679235063
transform 1 0 544 0 1 9484
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_6
timestamp 1679235063
transform 1 0 544 0 1 10069
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_7
timestamp 1679235063
transform -1 0 -27 0 -1 10102
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_8
timestamp 1679235063
transform -1 0 -27 0 1 9504
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_0
timestamp 1679235063
transform 1 0 110 0 1 6046
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_1
timestamp 1679235063
transform 1 0 544 0 1 9879
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_2
timestamp 1679235063
transform 1 0 544 0 1 10431
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_3
timestamp 1679235063
transform -1 0 -27 0 -1 10536
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180858  sky130_fd_pr__via_l1m1__example_5595914180858_4
timestamp 1679235063
transform -1 0 -27 0 1 9868
box 0 0 1 1
<< labels >>
flabel metal1 s 542 9482 654 9522 0 FreeSans 400 90 0 0 RB
port 2 nsew
flabel metal1 s 154 6046 188 6080 0 FreeSans 200 0 0 0 RA
port 1 nsew
<< properties >>
string GDS_END 3736600
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3733212
<< end >>
