magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -66 395 1122 897
rect -66 377 268 395
rect 777 377 1122 395
<< pwell >>
rect 304 317 715 335
rect 38 315 715 317
rect 38 283 788 315
rect 38 43 1052 283
rect -26 -43 1082 43
<< mvnmos >>
rect 117 207 217 291
rect 383 225 483 309
rect 539 225 639 309
rect 873 107 973 257
<< mvpmos >>
rect 131 463 231 613
rect 397 463 497 613
rect 553 463 653 613
rect 873 443 973 743
<< mvndiff >>
rect 330 297 383 309
rect 64 268 117 291
rect 64 234 72 268
rect 106 234 117 268
rect 64 207 117 234
rect 217 266 270 291
rect 217 232 228 266
rect 262 232 270 266
rect 217 207 270 232
rect 330 263 338 297
rect 372 263 383 297
rect 330 225 383 263
rect 483 267 539 309
rect 483 233 494 267
rect 528 233 539 267
rect 483 225 539 233
rect 639 289 689 309
rect 639 257 762 289
rect 639 241 873 257
rect 639 225 665 241
rect 657 207 665 225
rect 699 207 749 241
rect 783 207 828 241
rect 862 207 873 241
rect 657 173 873 207
rect 344 153 386 165
rect 344 119 352 153
rect 344 107 386 119
rect 657 139 665 173
rect 699 139 749 173
rect 783 139 828 173
rect 862 139 873 173
rect 657 107 873 139
rect 973 245 1026 257
rect 973 211 984 245
rect 1018 211 1026 245
rect 973 153 1026 211
rect 973 119 984 153
rect 1018 119 1026 153
rect 973 107 1026 119
<< mvpdiff >>
rect 156 731 198 743
rect 156 697 164 731
rect 156 685 198 697
rect 820 731 873 743
rect 820 697 828 731
rect 862 697 873 731
rect 820 657 873 697
rect 820 623 828 657
rect 862 623 873 657
rect 820 613 873 623
rect 78 601 131 613
rect 78 567 86 601
rect 120 567 131 601
rect 78 509 131 567
rect 78 475 86 509
rect 120 475 131 509
rect 78 463 131 475
rect 231 601 284 613
rect 231 567 242 601
rect 276 567 284 601
rect 231 509 284 567
rect 231 475 242 509
rect 276 475 284 509
rect 231 463 284 475
rect 344 597 397 613
rect 344 563 352 597
rect 386 563 397 597
rect 344 509 397 563
rect 344 475 352 509
rect 386 475 397 509
rect 344 463 397 475
rect 497 605 553 613
rect 497 571 508 605
rect 542 571 553 605
rect 497 507 553 571
rect 497 473 508 507
rect 542 473 553 507
rect 497 463 553 473
rect 653 605 873 613
rect 653 571 664 605
rect 698 571 748 605
rect 782 583 873 605
rect 782 571 828 583
rect 653 549 828 571
rect 862 549 873 583
rect 653 505 873 549
rect 653 471 664 505
rect 698 471 748 505
rect 782 471 828 505
rect 862 471 873 505
rect 653 463 873 471
rect 823 443 873 463
rect 973 727 1026 743
rect 973 693 984 727
rect 1018 693 1026 727
rect 973 652 1026 693
rect 973 618 984 652
rect 1018 618 1026 652
rect 973 571 1026 618
rect 973 537 984 571
rect 1018 537 1026 571
rect 973 491 1026 537
rect 973 457 984 491
rect 1018 457 1026 491
rect 973 443 1026 457
<< mvndiffc >>
rect 72 234 106 268
rect 228 232 262 266
rect 338 263 372 297
rect 494 233 528 267
rect 665 207 699 241
rect 749 207 783 241
rect 828 207 862 241
rect 352 119 386 153
rect 665 139 699 173
rect 749 139 783 173
rect 828 139 862 173
rect 984 211 1018 245
rect 984 119 1018 153
<< mvpdiffc >>
rect 164 697 198 731
rect 828 697 862 731
rect 828 623 862 657
rect 86 567 120 601
rect 86 475 120 509
rect 242 567 276 601
rect 242 475 276 509
rect 352 563 386 597
rect 352 475 386 509
rect 508 571 542 605
rect 508 473 542 507
rect 664 571 698 605
rect 748 571 782 605
rect 828 549 862 583
rect 664 471 698 505
rect 748 471 782 505
rect 828 471 862 505
rect 984 693 1018 727
rect 984 618 1018 652
rect 984 537 1018 571
rect 984 457 1018 491
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
<< poly >>
rect 873 743 973 769
rect 131 613 231 639
rect 397 613 497 639
rect 553 613 653 639
rect 131 397 231 463
rect 397 428 497 463
rect 553 428 653 463
rect 397 417 653 428
rect 397 405 639 417
rect 873 411 973 443
rect 131 381 327 397
rect 131 347 209 381
rect 243 347 277 381
rect 311 347 327 381
rect 131 329 327 347
rect 397 371 421 405
rect 455 371 489 405
rect 523 371 557 405
rect 591 371 639 405
rect 397 346 639 371
rect 383 345 639 346
rect 819 395 973 411
rect 819 361 836 395
rect 870 361 904 395
rect 938 361 973 395
rect 819 345 973 361
rect 131 319 217 329
rect 117 291 217 319
rect 383 309 483 345
rect 539 309 639 345
rect 873 257 973 345
rect 117 181 217 207
rect 383 199 483 225
rect 539 199 639 225
rect 873 77 973 107
<< polycont >>
rect 209 347 243 381
rect 277 347 311 381
rect 421 371 455 405
rect 489 371 523 405
rect 557 371 591 405
rect 836 361 870 395
rect 904 361 938 395
<< mvndiffres >>
rect 386 107 657 165
<< mvpdiffres >>
rect 198 685 820 743
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 148 731 206 747
rect 17 697 164 731
rect 198 697 206 731
rect 17 395 51 697
rect 148 681 206 697
rect 626 731 914 747
rect 626 729 828 731
rect 862 729 914 731
rect 626 695 645 729
rect 679 695 717 729
rect 751 695 789 729
rect 823 697 828 729
rect 823 695 861 697
rect 895 695 914 729
rect 626 681 914 695
rect 240 647 558 681
rect 86 601 136 617
rect 120 567 136 601
rect 86 509 136 567
rect 120 475 136 509
rect 86 467 136 475
rect 240 601 292 647
rect 240 567 242 601
rect 276 567 292 601
rect 240 509 292 567
rect 240 475 242 509
rect 276 475 292 509
rect 86 433 175 467
rect 240 459 292 475
rect 331 597 402 613
rect 331 563 352 597
rect 386 563 402 597
rect 331 509 402 563
rect 331 475 352 509
rect 386 475 402 509
rect 331 466 402 475
rect 492 605 558 647
rect 492 571 508 605
rect 542 571 558 605
rect 492 507 558 571
rect 492 473 508 507
rect 542 473 558 507
rect 17 361 106 395
rect 56 268 106 361
rect 56 234 72 268
rect 56 218 106 234
rect 141 159 175 433
rect 331 397 367 466
rect 492 464 558 473
rect 647 657 914 681
rect 647 623 828 657
rect 862 623 914 657
rect 647 605 914 623
rect 647 571 664 605
rect 698 571 748 605
rect 782 583 914 605
rect 782 571 828 583
rect 647 549 828 571
rect 862 549 914 583
rect 647 505 914 549
rect 647 471 664 505
rect 698 471 748 505
rect 782 471 828 505
rect 862 471 914 505
rect 647 464 914 471
rect 972 727 1039 743
rect 972 693 984 727
rect 1018 693 1039 727
rect 972 652 1039 693
rect 972 618 984 652
rect 1018 618 1039 652
rect 972 571 1039 618
rect 972 537 984 571
rect 1018 537 1039 571
rect 972 491 1039 537
rect 972 457 984 491
rect 1018 457 1039 491
rect 209 381 367 397
rect 243 347 277 381
rect 311 347 367 381
rect 403 405 661 430
rect 403 371 421 405
rect 455 371 489 405
rect 523 371 557 405
rect 591 371 661 405
rect 771 395 938 411
rect 209 337 367 347
rect 771 361 836 395
rect 870 361 904 395
rect 771 337 938 361
rect 209 331 938 337
rect 320 329 938 331
rect 320 301 842 329
rect 320 297 388 301
rect 212 266 278 282
rect 212 232 228 266
rect 262 232 278 266
rect 320 263 338 297
rect 372 263 388 297
rect 212 229 278 232
rect 478 233 494 267
rect 528 233 544 267
rect 478 229 544 233
rect 212 195 544 229
rect 624 241 926 257
rect 624 207 665 241
rect 699 207 749 241
rect 783 207 828 241
rect 862 207 926 241
rect 624 173 926 207
rect 141 153 402 159
rect 141 119 352 153
rect 386 119 402 153
rect 141 114 402 119
rect 624 139 665 173
rect 699 139 749 173
rect 783 139 828 173
rect 862 139 926 173
rect 624 119 926 139
rect 624 85 642 119
rect 676 85 714 119
rect 748 85 796 119
rect 830 85 882 119
rect 916 85 926 119
rect 972 245 1039 457
rect 972 211 984 245
rect 1018 211 1039 245
rect 972 153 1039 211
rect 972 119 984 153
rect 1018 119 1039 153
rect 972 103 1039 119
rect 624 75 926 85
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 645 695 679 729
rect 717 695 751 729
rect 789 695 823 729
rect 861 697 862 729
rect 862 697 895 729
rect 861 695 895 697
rect 642 85 676 119
rect 714 85 748 119
rect 796 85 830 119
rect 882 85 916 119
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 729 1056 763
rect 0 695 645 729
rect 679 695 717 729
rect 751 695 789 729
rect 823 695 861 729
rect 895 695 1056 729
rect 0 689 1056 695
rect 0 119 1056 125
rect 0 85 642 119
rect 676 85 714 119
rect 748 85 796 119
rect 830 85 882 119
rect 916 85 1056 119
rect 0 51 1056 85
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 schmittbuf_1
flabel comment s 121 718 121 718 0 FreeSans 200 0 0 0 resistive_li1_ok
flabel comment s 255 141 255 141 0 FreeSans 200 0 0 0 resistive_li1_ok
flabel locali s 991 168 1025 202 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 390 1025 424 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 464 1025 498 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 538 1025 572 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 991 612 1025 646 0 FreeSans 340 0 0 0 X
port 6 nsew signal output
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel metal1 s 0 689 1056 763 0 FreeSans 400 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 0 1056 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 791 1056 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel metal1 s 528 802 528 802 0 FreeSans 340 0 0 0 VPB
flabel metal1 s 0 51 1056 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 528 11 528 11 0 FreeSans 340 0 0 0 VNB
<< properties >>
string FIXED_BBOX 0 0 1056 814
string GDS_END 313324
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 301926
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
