magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< obsli1 >>
rect -3058 7901 3358 7983
rect -3058 -1900 -2976 7901
rect -1068 9 -934 5991
rect -830 9 -696 5991
rect 15 43 285 5957
rect 996 9 1130 5991
rect 1234 9 1368 5991
rect -209 -657 555 -443
rect 3276 -1900 3358 7901
rect -3058 -1982 3358 -1900
<< obsm1 >>
rect -3058 7901 3358 7983
rect -3058 -1900 -2976 7901
rect -1066 19 -936 5981
rect -828 19 -698 5981
rect 13 55 287 5945
rect 998 19 1128 5981
rect 1236 19 1366 5981
rect -209 -657 555 -443
rect 3276 -1900 3358 7901
rect -3058 -1982 3358 -1900
<< obsm2 >>
rect 22 57 278 5945
rect -209 -657 555 -443
<< properties >>
string FIXED_BBOX -3058 -1982 3358 7983
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8017720
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 7776368
<< end >>
