magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 94 21 367 157
rect 29 -17 63 17
<< locali >>
rect 31 326 75 487
rect 209 326 247 487
rect 31 292 351 326
rect 17 213 261 258
rect 295 179 351 292
rect 205 145 351 179
rect 205 56 250 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 109 459 175 493
rect 109 425 120 459
rect 154 425 175 459
rect 109 360 175 425
rect 281 459 347 493
rect 281 425 300 459
rect 334 425 347 459
rect 281 360 347 425
rect 112 17 171 122
rect 284 17 350 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 120 425 154 459
rect 300 425 334 459
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 14 459 354 468
rect 14 428 120 459
rect 108 425 120 428
rect 154 428 300 459
rect 154 425 166 428
rect 108 416 166 425
rect 288 425 300 428
rect 334 428 354 459
rect 334 425 346 428
rect 288 416 346 425
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
rlabel locali s 17 213 261 258 6 A
port 1 nsew signal input
rlabel metal1 s 288 416 346 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 108 416 166 428 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 14 428 354 468 6 KAPWR
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -48 368 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 205 56 250 145 6 Y
port 7 nsew signal output
rlabel locali s 205 145 351 179 6 Y
port 7 nsew signal output
rlabel locali s 295 179 351 292 6 Y
port 7 nsew signal output
rlabel locali s 31 292 351 326 6 Y
port 7 nsew signal output
rlabel locali s 209 326 247 487 6 Y
port 7 nsew signal output
rlabel locali s 31 326 75 487 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2285526
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2280822
<< end >>
