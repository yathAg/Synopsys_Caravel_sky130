magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect 0 0 564 1214
<< pmos >>
rect 204 102 254 1112
rect 310 102 360 1112
<< pdiff >>
rect 148 1100 204 1112
rect 148 1066 159 1100
rect 193 1066 204 1100
rect 148 1032 204 1066
rect 148 998 159 1032
rect 193 998 204 1032
rect 148 964 204 998
rect 148 930 159 964
rect 193 930 204 964
rect 148 896 204 930
rect 148 862 159 896
rect 193 862 204 896
rect 148 828 204 862
rect 148 794 159 828
rect 193 794 204 828
rect 148 760 204 794
rect 148 726 159 760
rect 193 726 204 760
rect 148 692 204 726
rect 148 658 159 692
rect 193 658 204 692
rect 148 624 204 658
rect 148 590 159 624
rect 193 590 204 624
rect 148 556 204 590
rect 148 522 159 556
rect 193 522 204 556
rect 148 488 204 522
rect 148 454 159 488
rect 193 454 204 488
rect 148 420 204 454
rect 148 386 159 420
rect 193 386 204 420
rect 148 352 204 386
rect 148 318 159 352
rect 193 318 204 352
rect 148 284 204 318
rect 148 250 159 284
rect 193 250 204 284
rect 148 216 204 250
rect 148 182 159 216
rect 193 182 204 216
rect 148 148 204 182
rect 148 114 159 148
rect 193 114 204 148
rect 148 102 204 114
rect 254 1100 310 1112
rect 254 1066 265 1100
rect 299 1066 310 1100
rect 254 1032 310 1066
rect 254 998 265 1032
rect 299 998 310 1032
rect 254 964 310 998
rect 254 930 265 964
rect 299 930 310 964
rect 254 896 310 930
rect 254 862 265 896
rect 299 862 310 896
rect 254 828 310 862
rect 254 794 265 828
rect 299 794 310 828
rect 254 760 310 794
rect 254 726 265 760
rect 299 726 310 760
rect 254 692 310 726
rect 254 658 265 692
rect 299 658 310 692
rect 254 624 310 658
rect 254 590 265 624
rect 299 590 310 624
rect 254 556 310 590
rect 254 522 265 556
rect 299 522 310 556
rect 254 488 310 522
rect 254 454 265 488
rect 299 454 310 488
rect 254 420 310 454
rect 254 386 265 420
rect 299 386 310 420
rect 254 352 310 386
rect 254 318 265 352
rect 299 318 310 352
rect 254 284 310 318
rect 254 250 265 284
rect 299 250 310 284
rect 254 216 310 250
rect 254 182 265 216
rect 299 182 310 216
rect 254 148 310 182
rect 254 114 265 148
rect 299 114 310 148
rect 254 102 310 114
rect 360 1100 416 1112
rect 360 1066 371 1100
rect 405 1066 416 1100
rect 360 1032 416 1066
rect 360 998 371 1032
rect 405 998 416 1032
rect 360 964 416 998
rect 360 930 371 964
rect 405 930 416 964
rect 360 896 416 930
rect 360 862 371 896
rect 405 862 416 896
rect 360 828 416 862
rect 360 794 371 828
rect 405 794 416 828
rect 360 760 416 794
rect 360 726 371 760
rect 405 726 416 760
rect 360 692 416 726
rect 360 658 371 692
rect 405 658 416 692
rect 360 624 416 658
rect 360 590 371 624
rect 405 590 416 624
rect 360 556 416 590
rect 360 522 371 556
rect 405 522 416 556
rect 360 488 416 522
rect 360 454 371 488
rect 405 454 416 488
rect 360 420 416 454
rect 360 386 371 420
rect 405 386 416 420
rect 360 352 416 386
rect 360 318 371 352
rect 405 318 416 352
rect 360 284 416 318
rect 360 250 371 284
rect 405 250 416 284
rect 360 216 416 250
rect 360 182 371 216
rect 405 182 416 216
rect 360 148 416 182
rect 360 114 371 148
rect 405 114 416 148
rect 360 102 416 114
<< pdiffc >>
rect 159 1066 193 1100
rect 159 998 193 1032
rect 159 930 193 964
rect 159 862 193 896
rect 159 794 193 828
rect 159 726 193 760
rect 159 658 193 692
rect 159 590 193 624
rect 159 522 193 556
rect 159 454 193 488
rect 159 386 193 420
rect 159 318 193 352
rect 159 250 193 284
rect 159 182 193 216
rect 159 114 193 148
rect 265 1066 299 1100
rect 265 998 299 1032
rect 265 930 299 964
rect 265 862 299 896
rect 265 794 299 828
rect 265 726 299 760
rect 265 658 299 692
rect 265 590 299 624
rect 265 522 299 556
rect 265 454 299 488
rect 265 386 299 420
rect 265 318 299 352
rect 265 250 299 284
rect 265 182 299 216
rect 265 114 299 148
rect 371 1066 405 1100
rect 371 998 405 1032
rect 371 930 405 964
rect 371 862 405 896
rect 371 794 405 828
rect 371 726 405 760
rect 371 658 405 692
rect 371 590 405 624
rect 371 522 405 556
rect 371 454 405 488
rect 371 386 405 420
rect 371 318 405 352
rect 371 250 405 284
rect 371 182 405 216
rect 371 114 405 148
<< nsubdiff >>
rect 36 1066 94 1112
rect 36 1032 48 1066
rect 82 1032 94 1066
rect 36 998 94 1032
rect 36 964 48 998
rect 82 964 94 998
rect 36 930 94 964
rect 36 896 48 930
rect 82 896 94 930
rect 36 862 94 896
rect 36 828 48 862
rect 82 828 94 862
rect 36 794 94 828
rect 36 760 48 794
rect 82 760 94 794
rect 36 726 94 760
rect 36 692 48 726
rect 82 692 94 726
rect 36 658 94 692
rect 36 624 48 658
rect 82 624 94 658
rect 36 590 94 624
rect 36 556 48 590
rect 82 556 94 590
rect 36 522 94 556
rect 36 488 48 522
rect 82 488 94 522
rect 36 454 94 488
rect 36 420 48 454
rect 82 420 94 454
rect 36 386 94 420
rect 36 352 48 386
rect 82 352 94 386
rect 36 318 94 352
rect 36 284 48 318
rect 82 284 94 318
rect 36 250 94 284
rect 36 216 48 250
rect 82 216 94 250
rect 36 182 94 216
rect 36 148 48 182
rect 82 148 94 182
rect 36 102 94 148
rect 470 1066 528 1112
rect 470 1032 482 1066
rect 516 1032 528 1066
rect 470 998 528 1032
rect 470 964 482 998
rect 516 964 528 998
rect 470 930 528 964
rect 470 896 482 930
rect 516 896 528 930
rect 470 862 528 896
rect 470 828 482 862
rect 516 828 528 862
rect 470 794 528 828
rect 470 760 482 794
rect 516 760 528 794
rect 470 726 528 760
rect 470 692 482 726
rect 516 692 528 726
rect 470 658 528 692
rect 470 624 482 658
rect 516 624 528 658
rect 470 590 528 624
rect 470 556 482 590
rect 516 556 528 590
rect 470 522 528 556
rect 470 488 482 522
rect 516 488 528 522
rect 470 454 528 488
rect 470 420 482 454
rect 516 420 528 454
rect 470 386 528 420
rect 470 352 482 386
rect 516 352 528 386
rect 470 318 528 352
rect 470 284 482 318
rect 516 284 528 318
rect 470 250 528 284
rect 470 216 482 250
rect 516 216 528 250
rect 470 182 528 216
rect 470 148 482 182
rect 516 148 528 182
rect 470 102 528 148
<< nsubdiffcont >>
rect 48 1032 82 1066
rect 48 964 82 998
rect 48 896 82 930
rect 48 828 82 862
rect 48 760 82 794
rect 48 692 82 726
rect 48 624 82 658
rect 48 556 82 590
rect 48 488 82 522
rect 48 420 82 454
rect 48 352 82 386
rect 48 284 82 318
rect 48 216 82 250
rect 48 148 82 182
rect 482 1032 516 1066
rect 482 964 516 998
rect 482 896 516 930
rect 482 828 516 862
rect 482 760 516 794
rect 482 692 516 726
rect 482 624 516 658
rect 482 556 516 590
rect 482 488 516 522
rect 482 420 516 454
rect 482 352 516 386
rect 482 284 516 318
rect 482 216 516 250
rect 482 148 516 182
<< poly >>
rect 181 1194 383 1214
rect 181 1160 197 1194
rect 231 1160 265 1194
rect 299 1160 333 1194
rect 367 1160 383 1194
rect 181 1144 383 1160
rect 204 1112 254 1144
rect 310 1112 360 1144
rect 204 70 254 102
rect 310 70 360 102
rect 181 54 383 70
rect 181 20 197 54
rect 231 20 265 54
rect 299 20 333 54
rect 367 20 383 54
rect 181 0 383 20
<< polycont >>
rect 197 1160 231 1194
rect 265 1160 299 1194
rect 333 1160 367 1194
rect 197 20 231 54
rect 265 20 299 54
rect 333 20 367 54
<< locali >>
rect 181 1160 193 1194
rect 231 1160 265 1194
rect 299 1160 333 1194
rect 371 1160 383 1194
rect 159 1100 193 1116
rect 48 1020 82 1032
rect 48 948 82 964
rect 48 876 82 896
rect 48 804 82 828
rect 48 732 82 760
rect 48 660 82 692
rect 48 590 82 624
rect 48 522 82 554
rect 48 454 82 482
rect 48 386 82 410
rect 48 318 82 338
rect 48 250 82 266
rect 48 182 82 194
rect 159 1032 193 1058
rect 159 964 193 986
rect 159 896 193 914
rect 159 828 193 842
rect 159 760 193 770
rect 159 692 193 698
rect 159 624 193 626
rect 159 588 193 590
rect 159 516 193 522
rect 159 444 193 454
rect 159 372 193 386
rect 159 300 193 318
rect 159 228 193 250
rect 159 156 193 182
rect 159 98 193 114
rect 265 1100 299 1116
rect 265 1032 299 1058
rect 265 964 299 986
rect 265 896 299 914
rect 265 828 299 842
rect 265 760 299 770
rect 265 692 299 698
rect 265 624 299 626
rect 265 588 299 590
rect 265 516 299 522
rect 265 444 299 454
rect 265 372 299 386
rect 265 300 299 318
rect 265 228 299 250
rect 265 156 299 182
rect 265 98 299 114
rect 371 1100 405 1116
rect 371 1032 405 1058
rect 371 964 405 986
rect 371 896 405 914
rect 371 828 405 842
rect 371 760 405 770
rect 371 692 405 698
rect 371 624 405 626
rect 371 588 405 590
rect 371 516 405 522
rect 371 444 405 454
rect 371 372 405 386
rect 371 300 405 318
rect 371 228 405 250
rect 371 156 405 182
rect 482 1020 516 1032
rect 482 948 516 964
rect 482 876 516 896
rect 482 804 516 828
rect 482 732 516 760
rect 482 660 516 692
rect 482 590 516 624
rect 482 522 516 554
rect 482 454 516 482
rect 482 386 516 410
rect 482 318 516 338
rect 482 250 516 266
rect 482 182 516 194
rect 371 98 405 114
rect 181 20 193 54
rect 231 20 265 54
rect 299 20 333 54
rect 371 20 383 54
<< viali >>
rect 193 1160 197 1194
rect 197 1160 227 1194
rect 265 1160 299 1194
rect 337 1160 367 1194
rect 367 1160 371 1194
rect 48 1066 82 1092
rect 48 1058 82 1066
rect 48 998 82 1020
rect 48 986 82 998
rect 48 930 82 948
rect 48 914 82 930
rect 48 862 82 876
rect 48 842 82 862
rect 48 794 82 804
rect 48 770 82 794
rect 48 726 82 732
rect 48 698 82 726
rect 48 658 82 660
rect 48 626 82 658
rect 48 556 82 588
rect 48 554 82 556
rect 48 488 82 516
rect 48 482 82 488
rect 48 420 82 444
rect 48 410 82 420
rect 48 352 82 372
rect 48 338 82 352
rect 48 284 82 300
rect 48 266 82 284
rect 48 216 82 228
rect 48 194 82 216
rect 48 148 82 156
rect 48 122 82 148
rect 159 1066 193 1092
rect 159 1058 193 1066
rect 159 998 193 1020
rect 159 986 193 998
rect 159 930 193 948
rect 159 914 193 930
rect 159 862 193 876
rect 159 842 193 862
rect 159 794 193 804
rect 159 770 193 794
rect 159 726 193 732
rect 159 698 193 726
rect 159 658 193 660
rect 159 626 193 658
rect 159 556 193 588
rect 159 554 193 556
rect 159 488 193 516
rect 159 482 193 488
rect 159 420 193 444
rect 159 410 193 420
rect 159 352 193 372
rect 159 338 193 352
rect 159 284 193 300
rect 159 266 193 284
rect 159 216 193 228
rect 159 194 193 216
rect 159 148 193 156
rect 159 122 193 148
rect 265 1066 299 1092
rect 265 1058 299 1066
rect 265 998 299 1020
rect 265 986 299 998
rect 265 930 299 948
rect 265 914 299 930
rect 265 862 299 876
rect 265 842 299 862
rect 265 794 299 804
rect 265 770 299 794
rect 265 726 299 732
rect 265 698 299 726
rect 265 658 299 660
rect 265 626 299 658
rect 265 556 299 588
rect 265 554 299 556
rect 265 488 299 516
rect 265 482 299 488
rect 265 420 299 444
rect 265 410 299 420
rect 265 352 299 372
rect 265 338 299 352
rect 265 284 299 300
rect 265 266 299 284
rect 265 216 299 228
rect 265 194 299 216
rect 265 148 299 156
rect 265 122 299 148
rect 371 1066 405 1092
rect 371 1058 405 1066
rect 371 998 405 1020
rect 371 986 405 998
rect 371 930 405 948
rect 371 914 405 930
rect 371 862 405 876
rect 371 842 405 862
rect 371 794 405 804
rect 371 770 405 794
rect 371 726 405 732
rect 371 698 405 726
rect 371 658 405 660
rect 371 626 405 658
rect 371 556 405 588
rect 371 554 405 556
rect 371 488 405 516
rect 371 482 405 488
rect 371 420 405 444
rect 371 410 405 420
rect 371 352 405 372
rect 371 338 405 352
rect 371 284 405 300
rect 371 266 405 284
rect 371 216 405 228
rect 371 194 405 216
rect 371 148 405 156
rect 371 122 405 148
rect 482 1066 516 1092
rect 482 1058 516 1066
rect 482 998 516 1020
rect 482 986 516 998
rect 482 930 516 948
rect 482 914 516 930
rect 482 862 516 876
rect 482 842 516 862
rect 482 794 516 804
rect 482 770 516 794
rect 482 726 516 732
rect 482 698 516 726
rect 482 658 516 660
rect 482 626 516 658
rect 482 556 516 588
rect 482 554 516 556
rect 482 488 516 516
rect 482 482 516 488
rect 482 420 516 444
rect 482 410 516 420
rect 482 352 516 372
rect 482 338 516 352
rect 482 284 516 300
rect 482 266 516 284
rect 482 216 516 228
rect 482 194 516 216
rect 482 148 516 156
rect 482 122 516 148
rect 193 20 197 54
rect 197 20 227 54
rect 265 20 299 54
rect 337 20 367 54
rect 367 20 371 54
<< metal1 >>
rect 181 1194 383 1214
rect 181 1160 193 1194
rect 227 1160 265 1194
rect 299 1160 337 1194
rect 371 1160 383 1194
rect 181 1148 383 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 156 94 194
rect 36 122 48 156
rect 82 122 94 156
rect 36 110 94 122
rect 150 1092 202 1104
rect 150 1058 159 1092
rect 193 1058 202 1092
rect 150 1020 202 1058
rect 150 986 159 1020
rect 193 986 202 1020
rect 150 948 202 986
rect 150 914 159 948
rect 193 914 202 948
rect 150 876 202 914
rect 150 842 159 876
rect 193 842 202 876
rect 150 804 202 842
rect 150 770 159 804
rect 193 770 202 804
rect 150 732 202 770
rect 150 698 159 732
rect 193 698 202 732
rect 150 660 202 698
rect 150 626 159 660
rect 193 626 202 660
rect 150 588 202 626
rect 150 554 159 588
rect 193 554 202 588
rect 150 552 202 554
rect 150 488 159 500
rect 193 488 202 500
rect 150 424 159 436
rect 193 424 202 436
rect 150 360 159 372
rect 193 360 202 372
rect 150 300 202 308
rect 150 296 159 300
rect 193 296 202 300
rect 150 232 202 244
rect 150 168 202 180
rect 150 110 202 116
rect 256 1098 308 1104
rect 256 1034 308 1046
rect 256 970 308 982
rect 256 914 265 918
rect 299 914 308 918
rect 256 906 308 914
rect 256 842 265 854
rect 299 842 308 854
rect 256 778 265 790
rect 299 778 308 790
rect 256 714 265 726
rect 299 714 308 726
rect 256 660 308 662
rect 256 626 265 660
rect 299 626 308 660
rect 256 588 308 626
rect 256 554 265 588
rect 299 554 308 588
rect 256 516 308 554
rect 256 482 265 516
rect 299 482 308 516
rect 256 444 308 482
rect 256 410 265 444
rect 299 410 308 444
rect 256 372 308 410
rect 256 338 265 372
rect 299 338 308 372
rect 256 300 308 338
rect 256 266 265 300
rect 299 266 308 300
rect 256 228 308 266
rect 256 194 265 228
rect 299 194 308 228
rect 256 156 308 194
rect 256 122 265 156
rect 299 122 308 156
rect 256 110 308 122
rect 362 1092 414 1104
rect 362 1058 371 1092
rect 405 1058 414 1092
rect 362 1020 414 1058
rect 362 986 371 1020
rect 405 986 414 1020
rect 362 948 414 986
rect 362 914 371 948
rect 405 914 414 948
rect 362 876 414 914
rect 362 842 371 876
rect 405 842 414 876
rect 362 804 414 842
rect 362 770 371 804
rect 405 770 414 804
rect 362 732 414 770
rect 362 698 371 732
rect 405 698 414 732
rect 362 660 414 698
rect 362 626 371 660
rect 405 626 414 660
rect 362 588 414 626
rect 362 554 371 588
rect 405 554 414 588
rect 362 552 414 554
rect 362 488 371 500
rect 405 488 414 500
rect 362 424 371 436
rect 405 424 414 436
rect 362 360 371 372
rect 405 360 414 372
rect 362 300 414 308
rect 362 296 371 300
rect 405 296 414 300
rect 362 232 414 244
rect 362 168 414 180
rect 362 110 414 116
rect 470 1092 528 1104
rect 470 1058 482 1092
rect 516 1058 528 1092
rect 470 1020 528 1058
rect 470 986 482 1020
rect 516 986 528 1020
rect 470 948 528 986
rect 470 914 482 948
rect 516 914 528 948
rect 470 876 528 914
rect 470 842 482 876
rect 516 842 528 876
rect 470 804 528 842
rect 470 770 482 804
rect 516 770 528 804
rect 470 732 528 770
rect 470 698 482 732
rect 516 698 528 732
rect 470 660 528 698
rect 470 626 482 660
rect 516 626 528 660
rect 470 588 528 626
rect 470 554 482 588
rect 516 554 528 588
rect 470 516 528 554
rect 470 482 482 516
rect 516 482 528 516
rect 470 444 528 482
rect 470 410 482 444
rect 516 410 528 444
rect 470 372 528 410
rect 470 338 482 372
rect 516 338 528 372
rect 470 300 528 338
rect 470 266 482 300
rect 516 266 528 300
rect 470 228 528 266
rect 470 194 482 228
rect 516 194 528 228
rect 470 156 528 194
rect 470 122 482 156
rect 516 122 528 156
rect 470 110 528 122
rect 181 54 383 66
rect 181 20 193 54
rect 227 20 265 54
rect 299 20 337 54
rect 371 20 383 54
rect 181 0 383 20
<< via1 >>
rect 150 516 202 552
rect 150 500 159 516
rect 159 500 193 516
rect 193 500 202 516
rect 150 482 159 488
rect 159 482 193 488
rect 193 482 202 488
rect 150 444 202 482
rect 150 436 159 444
rect 159 436 193 444
rect 193 436 202 444
rect 150 410 159 424
rect 159 410 193 424
rect 193 410 202 424
rect 150 372 202 410
rect 150 338 159 360
rect 159 338 193 360
rect 193 338 202 360
rect 150 308 202 338
rect 150 266 159 296
rect 159 266 193 296
rect 193 266 202 296
rect 150 244 202 266
rect 150 228 202 232
rect 150 194 159 228
rect 159 194 193 228
rect 193 194 202 228
rect 150 180 202 194
rect 150 156 202 168
rect 150 122 159 156
rect 159 122 193 156
rect 193 122 202 156
rect 150 116 202 122
rect 256 1092 308 1098
rect 256 1058 265 1092
rect 265 1058 299 1092
rect 299 1058 308 1092
rect 256 1046 308 1058
rect 256 1020 308 1034
rect 256 986 265 1020
rect 265 986 299 1020
rect 299 986 308 1020
rect 256 982 308 986
rect 256 948 308 970
rect 256 918 265 948
rect 265 918 299 948
rect 299 918 308 948
rect 256 876 308 906
rect 256 854 265 876
rect 265 854 299 876
rect 299 854 308 876
rect 256 804 308 842
rect 256 790 265 804
rect 265 790 299 804
rect 299 790 308 804
rect 256 770 265 778
rect 265 770 299 778
rect 299 770 308 778
rect 256 732 308 770
rect 256 726 265 732
rect 265 726 299 732
rect 299 726 308 732
rect 256 698 265 714
rect 265 698 299 714
rect 299 698 308 714
rect 256 662 308 698
rect 362 516 414 552
rect 362 500 371 516
rect 371 500 405 516
rect 405 500 414 516
rect 362 482 371 488
rect 371 482 405 488
rect 405 482 414 488
rect 362 444 414 482
rect 362 436 371 444
rect 371 436 405 444
rect 405 436 414 444
rect 362 410 371 424
rect 371 410 405 424
rect 405 410 414 424
rect 362 372 414 410
rect 362 338 371 360
rect 371 338 405 360
rect 405 338 414 360
rect 362 308 414 338
rect 362 266 371 296
rect 371 266 405 296
rect 405 266 414 296
rect 362 244 414 266
rect 362 228 414 232
rect 362 194 371 228
rect 371 194 405 228
rect 405 194 414 228
rect 362 180 414 194
rect 362 156 414 168
rect 362 122 371 156
rect 371 122 405 156
rect 405 122 414 156
rect 362 116 414 122
<< metal2 >>
rect 10 1098 554 1104
rect 10 1046 256 1098
rect 308 1046 554 1098
rect 10 1034 554 1046
rect 10 982 256 1034
rect 308 982 554 1034
rect 10 970 554 982
rect 10 918 256 970
rect 308 918 554 970
rect 10 906 554 918
rect 10 854 256 906
rect 308 854 554 906
rect 10 842 554 854
rect 10 790 256 842
rect 308 790 554 842
rect 10 778 554 790
rect 10 726 256 778
rect 308 726 554 778
rect 10 714 554 726
rect 10 662 256 714
rect 308 662 554 714
rect 10 632 554 662
rect 10 552 554 582
rect 10 500 150 552
rect 202 500 362 552
rect 414 500 554 552
rect 10 488 554 500
rect 10 436 150 488
rect 202 436 362 488
rect 414 436 554 488
rect 10 424 554 436
rect 10 372 150 424
rect 202 372 362 424
rect 414 372 554 424
rect 10 360 554 372
rect 10 308 150 360
rect 202 308 362 360
rect 414 308 554 360
rect 10 296 554 308
rect 10 244 150 296
rect 202 244 362 296
rect 414 244 554 296
rect 10 232 554 244
rect 10 180 150 232
rect 202 180 362 232
rect 414 180 554 232
rect 10 168 554 180
rect 10 116 150 168
rect 202 116 362 168
rect 414 116 554 168
rect 10 110 554 116
<< labels >>
flabel metal2 s 16 317 37 381 0 FreeSans 400 90 0 0 SOURCE
port 2 nsew
flabel metal2 s 15 799 34 869 0 FreeSans 400 90 0 0 DRAIN
port 3 nsew
flabel metal1 s 181 1148 383 1214 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 181 0 383 66 0 FreeSans 300 0 0 0 GATE
port 4 nsew
flabel metal1 s 496 732 496 732 7 FreeSans 400 90 0 0 BULK
flabel metal1 s 60 732 60 732 7 FreeSans 400 90 0 0 BULK
<< properties >>
string GDS_END 9331582
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9316058
<< end >>
