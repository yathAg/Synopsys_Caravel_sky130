magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 366 157 827 203
rect 1 21 827 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 184 47 214 131
rect 444 47 474 177
rect 528 47 558 177
rect 635 47 665 177
rect 719 47 749 177
<< scpmoshvt >>
rect 79 369 109 497
rect 184 369 214 497
rect 372 309 402 497
rect 456 309 486 497
rect 635 297 665 497
rect 719 297 749 497
<< ndiff >>
rect 27 106 79 131
rect 27 72 35 106
rect 69 72 79 106
rect 27 47 79 72
rect 109 89 184 131
rect 109 55 119 89
rect 153 55 184 89
rect 109 47 184 55
rect 214 106 266 131
rect 214 72 224 106
rect 258 72 266 106
rect 214 47 266 72
rect 392 129 444 177
rect 392 95 400 129
rect 434 95 444 129
rect 392 47 444 95
rect 474 89 528 177
rect 474 55 484 89
rect 518 55 528 89
rect 474 47 528 55
rect 558 129 635 177
rect 558 95 579 129
rect 613 95 635 129
rect 558 47 635 95
rect 665 169 719 177
rect 665 135 675 169
rect 709 135 719 169
rect 665 47 719 135
rect 749 93 801 177
rect 749 59 759 93
rect 793 59 801 93
rect 749 47 801 59
<< pdiff >>
rect 27 461 79 497
rect 27 427 35 461
rect 69 427 79 461
rect 27 369 79 427
rect 109 489 184 497
rect 109 455 130 489
rect 164 455 184 489
rect 109 421 184 455
rect 109 387 130 421
rect 164 387 184 421
rect 109 369 184 387
rect 214 461 266 497
rect 214 427 224 461
rect 258 427 266 461
rect 214 369 266 427
rect 320 477 372 497
rect 320 443 328 477
rect 362 443 372 477
rect 320 309 372 443
rect 402 489 456 497
rect 402 455 412 489
rect 446 455 456 489
rect 402 309 456 455
rect 486 477 635 497
rect 486 443 508 477
rect 542 443 576 477
rect 610 443 635 477
rect 486 309 635 443
rect 501 297 635 309
rect 665 416 719 497
rect 665 382 675 416
rect 709 382 719 416
rect 665 348 719 382
rect 665 314 675 348
rect 709 314 719 348
rect 665 297 719 314
rect 749 477 801 497
rect 749 443 759 477
rect 793 443 801 477
rect 749 409 801 443
rect 749 375 759 409
rect 793 375 801 409
rect 749 297 801 375
<< ndiffc >>
rect 35 72 69 106
rect 119 55 153 89
rect 224 72 258 106
rect 400 95 434 129
rect 484 55 518 89
rect 579 95 613 129
rect 675 135 709 169
rect 759 59 793 93
<< pdiffc >>
rect 35 427 69 461
rect 130 455 164 489
rect 130 387 164 421
rect 224 427 258 461
rect 328 443 362 477
rect 412 455 446 489
rect 508 443 542 477
rect 576 443 610 477
rect 675 382 709 416
rect 675 314 709 348
rect 759 443 793 477
rect 759 375 793 409
<< poly >>
rect 79 497 109 523
rect 184 497 214 523
rect 372 497 402 523
rect 456 497 486 523
rect 635 497 665 523
rect 719 497 749 523
rect 79 265 109 369
rect 184 294 214 369
rect 372 294 402 309
rect 456 294 486 309
rect 184 272 486 294
rect 79 249 142 265
rect 79 215 98 249
rect 132 215 142 249
rect 79 199 142 215
rect 184 264 485 272
rect 184 249 256 264
rect 635 259 665 297
rect 719 259 749 297
rect 184 215 206 249
rect 240 215 256 249
rect 527 249 593 259
rect 527 222 543 249
rect 184 205 256 215
rect 444 215 543 222
rect 577 215 593 249
rect 79 131 109 199
rect 184 131 214 205
rect 444 192 593 215
rect 635 249 749 259
rect 635 215 675 249
rect 709 215 749 249
rect 635 205 749 215
rect 444 177 474 192
rect 528 177 558 192
rect 635 177 665 205
rect 719 177 749 205
rect 79 21 109 47
rect 184 21 214 47
rect 444 21 474 47
rect 528 21 558 47
rect 635 21 665 47
rect 719 21 749 47
<< polycont >>
rect 98 215 132 249
rect 206 215 240 249
rect 543 215 577 249
rect 675 215 709 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 461 69 493
rect 17 427 35 461
rect 17 369 69 427
rect 103 489 190 527
rect 103 455 130 489
rect 164 455 190 489
rect 103 421 190 455
rect 103 387 130 421
rect 164 387 190 421
rect 103 369 190 387
rect 224 461 282 493
rect 258 427 282 461
rect 17 255 64 369
rect 224 353 282 427
rect 320 477 362 493
rect 320 443 328 477
rect 396 489 462 527
rect 396 455 412 489
rect 446 455 462 489
rect 496 477 811 493
rect 320 421 362 443
rect 496 443 508 477
rect 542 443 576 477
rect 610 459 759 477
rect 610 443 625 459
rect 496 421 625 443
rect 793 443 811 477
rect 320 387 625 421
rect 659 416 725 425
rect 659 382 675 416
rect 709 382 725 416
rect 659 353 725 382
rect 759 409 811 443
rect 793 375 811 409
rect 759 359 811 375
rect 17 221 30 255
rect 17 123 64 221
rect 98 249 156 335
rect 224 289 347 353
rect 381 348 725 353
rect 381 314 675 348
rect 709 325 725 348
rect 709 314 811 325
rect 381 289 811 314
rect 290 255 347 289
rect 132 215 156 249
rect 98 153 156 215
rect 190 249 256 255
rect 190 215 206 249
rect 240 215 256 249
rect 190 153 256 215
rect 290 249 593 255
rect 290 215 543 249
rect 577 215 593 249
rect 290 205 593 215
rect 649 249 676 255
rect 649 215 675 249
rect 710 221 731 255
rect 709 215 731 221
rect 649 205 731 215
rect 17 106 69 123
rect 290 119 346 205
rect 765 171 811 289
rect 17 72 35 106
rect 17 56 69 72
rect 103 89 170 119
rect 103 55 119 89
rect 153 55 170 89
rect 103 17 170 55
rect 204 106 346 119
rect 204 72 224 106
rect 258 72 346 106
rect 204 51 346 72
rect 380 131 625 171
rect 380 129 434 131
rect 380 95 400 129
rect 568 129 625 131
rect 380 51 434 95
rect 468 89 534 97
rect 468 55 484 89
rect 518 55 534 89
rect 568 95 579 129
rect 613 95 625 129
rect 659 169 811 171
rect 659 135 675 169
rect 709 135 811 169
rect 659 127 811 135
rect 568 93 625 95
rect 568 59 759 93
rect 793 59 810 93
rect 568 55 810 59
rect 468 17 534 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 30 221 64 255
rect 676 249 710 255
rect 676 221 709 249
rect 709 221 710 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 17 255 76 261
rect 17 221 30 255
rect 64 252 76 255
rect 664 255 722 261
rect 664 252 676 255
rect 64 224 676 252
rect 64 221 76 224
rect 17 215 76 221
rect 664 221 676 224
rect 710 221 722 255
rect 664 215 722 221
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 768 221 802 255 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 768 289 802 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 122 153 156 187 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 676 357 710 391 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 122 289 156 323 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 TE_B
port 2 nsew signal input
flabel locali s 584 289 618 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 493 289 526 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 402 289 436 323 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel locali s 768 153 802 187 0 FreeSans 200 0 0 0 Z
port 7 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 4 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 5 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 3 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 6 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 ebufn_2
rlabel metal1 s 0 -48 828 48 1 VGND
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 6 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 2946808
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2939612
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
