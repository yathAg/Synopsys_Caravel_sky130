magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< pwell >>
rect 15 163 811 545
<< nmos >>
rect 171 189 201 519
rect 257 189 293 519
rect 349 189 385 519
rect 441 189 477 519
rect 533 189 569 519
rect 625 189 655 519
<< ndiff >>
rect 111 507 171 519
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 507 257 519
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 293 507 349 519
rect 293 473 304 507
rect 338 473 349 507
rect 293 439 349 473
rect 293 405 304 439
rect 338 405 349 439
rect 293 371 349 405
rect 293 337 304 371
rect 338 337 349 371
rect 293 303 349 337
rect 293 269 304 303
rect 338 269 349 303
rect 293 235 349 269
rect 293 201 304 235
rect 338 201 349 235
rect 293 189 349 201
rect 385 507 441 519
rect 385 473 396 507
rect 430 473 441 507
rect 385 439 441 473
rect 385 405 396 439
rect 430 405 441 439
rect 385 371 441 405
rect 385 337 396 371
rect 430 337 441 371
rect 385 303 441 337
rect 385 269 396 303
rect 430 269 441 303
rect 385 235 441 269
rect 385 201 396 235
rect 430 201 441 235
rect 385 189 441 201
rect 477 507 533 519
rect 477 473 488 507
rect 522 473 533 507
rect 477 439 533 473
rect 477 405 488 439
rect 522 405 533 439
rect 477 371 533 405
rect 477 337 488 371
rect 522 337 533 371
rect 477 303 533 337
rect 477 269 488 303
rect 522 269 533 303
rect 477 235 533 269
rect 477 201 488 235
rect 522 201 533 235
rect 477 189 533 201
rect 569 507 625 519
rect 569 473 580 507
rect 614 473 625 507
rect 569 439 625 473
rect 569 405 580 439
rect 614 405 625 439
rect 569 371 625 405
rect 569 337 580 371
rect 614 337 625 371
rect 569 303 625 337
rect 569 269 580 303
rect 614 269 625 303
rect 569 235 625 269
rect 569 201 580 235
rect 614 201 625 235
rect 569 189 625 201
rect 655 507 715 519
rect 655 473 666 507
rect 700 473 715 507
rect 655 439 715 473
rect 655 405 666 439
rect 700 405 715 439
rect 655 371 715 405
rect 655 337 666 371
rect 700 337 715 371
rect 655 303 715 337
rect 655 269 666 303
rect 700 269 715 303
rect 655 235 715 269
rect 655 201 666 235
rect 700 201 715 235
rect 655 189 715 201
<< ndiffc >>
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 304 473 338 507
rect 304 405 338 439
rect 304 337 338 371
rect 304 269 338 303
rect 304 201 338 235
rect 396 473 430 507
rect 396 405 430 439
rect 396 337 430 371
rect 396 269 430 303
rect 396 201 430 235
rect 488 473 522 507
rect 488 405 522 439
rect 488 337 522 371
rect 488 269 522 303
rect 488 201 522 235
rect 580 473 614 507
rect 580 405 614 439
rect 580 337 614 371
rect 580 269 614 303
rect 580 201 614 235
rect 666 473 700 507
rect 666 405 700 439
rect 666 337 700 371
rect 666 269 700 303
rect 666 201 700 235
<< psubdiff >>
rect 41 507 111 519
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 715 507 785 519
rect 715 473 734 507
rect 768 473 785 507
rect 715 439 785 473
rect 715 405 734 439
rect 768 405 785 439
rect 715 371 785 405
rect 715 337 734 371
rect 768 337 785 371
rect 715 303 785 337
rect 715 269 734 303
rect 768 269 785 303
rect 715 235 785 269
rect 715 201 734 235
rect 768 201 785 235
rect 715 189 785 201
<< psubdiffcont >>
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 734 473 768 507
rect 734 405 768 439
rect 734 337 768 371
rect 734 269 768 303
rect 734 201 768 235
<< poly >>
rect 243 687 583 708
rect 116 595 201 611
rect 116 561 132 595
rect 166 561 201 595
rect 243 585 260 687
rect 566 585 583 687
rect 243 569 583 585
rect 625 595 710 611
rect 116 545 201 561
rect 171 519 201 545
rect 257 519 293 569
rect 349 519 385 569
rect 441 519 477 569
rect 533 519 569 569
rect 625 561 660 595
rect 694 561 710 595
rect 625 545 710 561
rect 625 519 655 545
rect 171 163 201 189
rect 116 147 201 163
rect 116 113 132 147
rect 166 113 201 147
rect 257 139 293 189
rect 349 139 385 189
rect 441 139 477 189
rect 533 139 569 189
rect 625 163 655 189
rect 625 147 710 163
rect 116 97 201 113
rect 243 123 583 139
rect 243 21 260 123
rect 566 21 583 123
rect 625 113 660 147
rect 694 113 710 147
rect 625 97 710 113
rect 243 0 583 21
<< polycont >>
rect 132 561 166 595
rect 260 585 566 687
rect 660 561 694 595
rect 132 113 166 147
rect 260 21 566 123
rect 660 113 694 147
<< locali >>
rect 238 689 588 708
rect 116 595 182 611
rect 116 561 132 595
rect 166 561 182 595
rect 238 583 252 689
rect 574 583 588 689
rect 238 569 588 583
rect 644 595 710 611
rect 116 545 182 561
rect 644 561 660 595
rect 694 561 710 595
rect 644 545 710 561
rect 116 523 160 545
rect 666 523 710 545
rect 41 507 160 523
rect 41 473 58 507
rect 92 479 126 507
rect 94 473 126 479
rect 41 445 60 473
rect 94 445 160 473
rect 41 439 160 445
rect 41 405 58 439
rect 92 407 126 439
rect 94 405 126 407
rect 41 373 60 405
rect 94 373 160 405
rect 41 371 160 373
rect 41 337 58 371
rect 92 337 126 371
rect 41 335 160 337
rect 41 303 60 335
rect 94 303 160 335
rect 41 269 58 303
rect 94 301 126 303
rect 92 269 126 301
rect 41 263 160 269
rect 41 235 60 263
rect 94 235 160 263
rect 41 201 58 235
rect 94 229 126 235
rect 92 201 126 229
rect 41 185 160 201
rect 212 507 246 523
rect 212 439 246 445
rect 212 371 246 373
rect 212 335 246 337
rect 212 263 246 269
rect 212 185 246 201
rect 304 507 338 523
rect 304 439 338 445
rect 304 371 338 373
rect 304 335 338 337
rect 304 263 338 269
rect 304 185 338 201
rect 396 507 430 523
rect 396 439 430 445
rect 396 371 430 373
rect 396 335 430 337
rect 396 263 430 269
rect 396 185 430 201
rect 488 507 522 523
rect 488 439 522 445
rect 488 371 522 373
rect 488 335 522 337
rect 488 263 522 269
rect 488 185 522 201
rect 580 507 614 523
rect 580 439 614 445
rect 580 371 614 373
rect 580 335 614 337
rect 580 263 614 269
rect 580 185 614 201
rect 666 507 785 523
rect 700 479 734 507
rect 700 473 732 479
rect 768 473 785 507
rect 666 445 732 473
rect 766 445 785 473
rect 666 439 785 445
rect 700 407 734 439
rect 700 405 732 407
rect 768 405 785 439
rect 666 373 732 405
rect 766 373 785 405
rect 666 371 785 373
rect 700 337 734 371
rect 768 337 785 371
rect 666 335 785 337
rect 666 303 732 335
rect 766 303 785 335
rect 700 301 732 303
rect 700 269 734 301
rect 768 269 785 303
rect 666 263 785 269
rect 666 235 732 263
rect 766 235 785 263
rect 700 229 732 235
rect 700 201 734 229
rect 768 201 785 235
rect 666 185 785 201
rect 116 163 160 185
rect 666 163 710 185
rect 116 147 182 163
rect 116 113 132 147
rect 166 113 182 147
rect 644 147 710 163
rect 116 97 182 113
rect 238 125 588 139
rect 238 19 252 125
rect 574 19 588 125
rect 644 113 660 147
rect 694 113 710 147
rect 644 97 710 113
rect 238 0 588 19
<< viali >>
rect 252 687 574 689
rect 252 585 260 687
rect 260 585 566 687
rect 566 585 574 687
rect 252 583 574 585
rect 60 473 92 479
rect 92 473 94 479
rect 60 445 94 473
rect 60 405 92 407
rect 92 405 94 407
rect 60 373 94 405
rect 60 303 94 335
rect 60 301 92 303
rect 92 301 94 303
rect 60 235 94 263
rect 60 229 92 235
rect 92 229 94 235
rect 212 473 246 479
rect 212 445 246 473
rect 212 405 246 407
rect 212 373 246 405
rect 212 303 246 335
rect 212 301 246 303
rect 212 235 246 263
rect 212 229 246 235
rect 304 473 338 479
rect 304 445 338 473
rect 304 405 338 407
rect 304 373 338 405
rect 304 303 338 335
rect 304 301 338 303
rect 304 235 338 263
rect 304 229 338 235
rect 396 473 430 479
rect 396 445 430 473
rect 396 405 430 407
rect 396 373 430 405
rect 396 303 430 335
rect 396 301 430 303
rect 396 235 430 263
rect 396 229 430 235
rect 488 473 522 479
rect 488 445 522 473
rect 488 405 522 407
rect 488 373 522 405
rect 488 303 522 335
rect 488 301 522 303
rect 488 235 522 263
rect 488 229 522 235
rect 580 473 614 479
rect 580 445 614 473
rect 580 405 614 407
rect 580 373 614 405
rect 580 303 614 335
rect 580 301 614 303
rect 580 235 614 263
rect 580 229 614 235
rect 732 473 734 479
rect 734 473 766 479
rect 732 445 766 473
rect 732 405 734 407
rect 734 405 766 407
rect 732 373 766 405
rect 732 303 766 335
rect 732 301 734 303
rect 734 301 766 303
rect 732 235 766 263
rect 732 229 734 235
rect 734 229 766 235
rect 252 123 574 125
rect 252 21 260 123
rect 260 21 566 123
rect 566 21 574 123
rect 252 19 574 21
<< metal1 >>
rect 236 689 590 708
rect 236 583 252 689
rect 574 583 590 689
rect 236 571 590 583
rect 41 479 100 507
rect 41 445 60 479
rect 94 445 100 479
rect 41 407 100 445
rect 41 373 60 407
rect 94 373 100 407
rect 41 335 100 373
rect 41 301 60 335
rect 94 301 100 335
rect 41 263 100 301
rect 41 229 60 263
rect 94 229 100 263
rect 41 201 100 229
rect 203 479 255 507
rect 203 445 212 479
rect 246 445 255 479
rect 203 407 255 445
rect 203 373 212 407
rect 246 373 255 407
rect 203 335 255 373
rect 203 323 212 335
rect 246 323 255 335
rect 203 263 255 271
rect 203 259 212 263
rect 246 259 255 263
rect 203 201 255 207
rect 295 501 347 507
rect 295 445 304 449
rect 338 445 347 449
rect 295 437 347 445
rect 295 373 304 385
rect 338 373 347 385
rect 295 335 347 373
rect 295 301 304 335
rect 338 301 347 335
rect 295 263 347 301
rect 295 229 304 263
rect 338 229 347 263
rect 295 201 347 229
rect 387 479 439 507
rect 387 445 396 479
rect 430 445 439 479
rect 387 407 439 445
rect 387 373 396 407
rect 430 373 439 407
rect 387 335 439 373
rect 387 323 396 335
rect 430 323 439 335
rect 387 263 439 271
rect 387 259 396 263
rect 430 259 439 263
rect 387 201 439 207
rect 479 501 531 507
rect 479 445 488 449
rect 522 445 531 449
rect 479 437 531 445
rect 479 373 488 385
rect 522 373 531 385
rect 479 335 531 373
rect 479 301 488 335
rect 522 301 531 335
rect 479 263 531 301
rect 479 229 488 263
rect 522 229 531 263
rect 479 201 531 229
rect 571 479 623 507
rect 571 445 580 479
rect 614 445 623 479
rect 571 407 623 445
rect 571 373 580 407
rect 614 373 623 407
rect 571 335 623 373
rect 571 323 580 335
rect 614 323 623 335
rect 571 263 623 271
rect 571 259 580 263
rect 614 259 623 263
rect 571 201 623 207
rect 726 479 785 507
rect 726 445 732 479
rect 766 445 785 479
rect 726 407 785 445
rect 726 373 732 407
rect 766 373 785 407
rect 726 335 785 373
rect 726 301 732 335
rect 766 301 785 335
rect 726 263 785 301
rect 726 229 732 263
rect 766 229 785 263
rect 726 201 785 229
rect 236 125 590 137
rect 236 19 252 125
rect 574 19 590 125
rect 236 0 590 19
<< via1 >>
rect 203 301 212 323
rect 212 301 246 323
rect 246 301 255 323
rect 203 271 255 301
rect 203 229 212 259
rect 212 229 246 259
rect 246 229 255 259
rect 203 207 255 229
rect 295 479 347 501
rect 295 449 304 479
rect 304 449 338 479
rect 338 449 347 479
rect 295 407 347 437
rect 295 385 304 407
rect 304 385 338 407
rect 338 385 347 407
rect 387 301 396 323
rect 396 301 430 323
rect 430 301 439 323
rect 387 271 439 301
rect 387 229 396 259
rect 396 229 430 259
rect 430 229 439 259
rect 387 207 439 229
rect 479 479 531 501
rect 479 449 488 479
rect 488 449 522 479
rect 522 449 531 479
rect 479 407 531 437
rect 479 385 488 407
rect 488 385 522 407
rect 522 385 531 407
rect 571 301 580 323
rect 580 301 614 323
rect 614 301 623 323
rect 571 271 623 301
rect 571 229 580 259
rect 580 229 614 259
rect 614 229 623 259
rect 571 207 623 229
<< metal2 >>
rect 14 501 812 507
rect 14 449 295 501
rect 347 449 479 501
rect 531 449 812 501
rect 14 437 812 449
rect 14 385 295 437
rect 347 385 479 437
rect 531 385 812 437
rect 14 379 812 385
rect 14 323 812 329
rect 14 271 203 323
rect 255 271 387 323
rect 439 271 571 323
rect 623 271 812 323
rect 14 259 812 271
rect 14 207 203 259
rect 255 207 387 259
rect 439 207 571 259
rect 623 207 812 259
rect 14 201 812 207
<< labels >>
flabel comment s 183 335 183 335 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 636 321 636 321 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 301 606 535 656 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 301 42 535 92 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 339 87 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 739 339 785 369 0 FreeSans 200 90 0 0 SUBSTRATE
port 4 nsew
flabel metal2 s 14 201 35 329 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 379 35 507 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 5725752
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 5710380
string device primitive
<< end >>
