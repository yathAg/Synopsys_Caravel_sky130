magic
tech sky130A
timestamp 1679235063
<< properties >>
string GDS_END 27764764
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27764504
<< end >>
