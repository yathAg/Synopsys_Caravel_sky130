magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< dnwell >>
rect 214 214 1978 3178
<< nwell >>
rect 134 2898 2058 3258
rect 134 494 494 2898
rect 1698 494 2058 2898
rect 134 134 2058 494
<< pwell >>
rect 0 3258 2192 3392
rect 0 134 134 3258
rect 628 628 1564 2764
rect 2058 134 2192 3258
rect 0 0 2192 134
<< ndiff >>
rect 896 2461 1296 2496
rect 896 931 909 2461
rect 1283 931 1296 2461
rect 896 896 1296 931
<< ndiffc >>
rect 909 931 1283 2461
<< psubdiff >>
rect 26 3342 2166 3366
rect 26 3308 50 3342
rect 84 3308 127 3342
rect 161 3308 195 3342
rect 229 3308 263 3342
rect 297 3308 331 3342
rect 365 3308 399 3342
rect 433 3308 467 3342
rect 501 3308 535 3342
rect 569 3308 603 3342
rect 637 3308 671 3342
rect 705 3308 739 3342
rect 773 3308 807 3342
rect 841 3308 875 3342
rect 909 3308 943 3342
rect 977 3308 1011 3342
rect 1045 3308 1079 3342
rect 1113 3308 1147 3342
rect 1181 3308 1215 3342
rect 1249 3308 1283 3342
rect 1317 3308 1351 3342
rect 1385 3308 1419 3342
rect 1453 3308 1487 3342
rect 1521 3308 1555 3342
rect 1589 3308 1623 3342
rect 1657 3308 1691 3342
rect 1725 3308 1759 3342
rect 1793 3308 1827 3342
rect 1861 3308 1895 3342
rect 1929 3308 1963 3342
rect 1997 3308 2031 3342
rect 2065 3308 2108 3342
rect 2142 3308 2166 3342
rect 26 3284 2166 3308
rect 26 3243 108 3284
rect 26 3209 50 3243
rect 84 3209 108 3243
rect 26 3175 108 3209
rect 26 3141 50 3175
rect 84 3141 108 3175
rect 26 3107 108 3141
rect 2084 3243 2166 3284
rect 2084 3209 2108 3243
rect 2142 3209 2166 3243
rect 2084 3175 2166 3209
rect 2084 3141 2108 3175
rect 2142 3141 2166 3175
rect 26 3073 50 3107
rect 84 3073 108 3107
rect 26 3039 108 3073
rect 26 3005 50 3039
rect 84 3005 108 3039
rect 26 2971 108 3005
rect 26 2937 50 2971
rect 84 2937 108 2971
rect 26 2903 108 2937
rect 26 2869 50 2903
rect 84 2869 108 2903
rect 26 2835 108 2869
rect 26 2801 50 2835
rect 84 2801 108 2835
rect 26 2767 108 2801
rect 26 2733 50 2767
rect 84 2733 108 2767
rect 26 2699 108 2733
rect 26 2665 50 2699
rect 84 2665 108 2699
rect 26 2631 108 2665
rect 26 2597 50 2631
rect 84 2597 108 2631
rect 26 2563 108 2597
rect 26 2529 50 2563
rect 84 2529 108 2563
rect 26 2495 108 2529
rect 26 2461 50 2495
rect 84 2461 108 2495
rect 26 2427 108 2461
rect 26 2393 50 2427
rect 84 2393 108 2427
rect 26 2359 108 2393
rect 26 2325 50 2359
rect 84 2325 108 2359
rect 26 2291 108 2325
rect 26 2257 50 2291
rect 84 2257 108 2291
rect 26 2223 108 2257
rect 26 2189 50 2223
rect 84 2189 108 2223
rect 26 2155 108 2189
rect 26 2121 50 2155
rect 84 2121 108 2155
rect 26 2087 108 2121
rect 26 2053 50 2087
rect 84 2053 108 2087
rect 26 2019 108 2053
rect 26 1985 50 2019
rect 84 1985 108 2019
rect 26 1951 108 1985
rect 26 1917 50 1951
rect 84 1917 108 1951
rect 26 1883 108 1917
rect 26 1849 50 1883
rect 84 1849 108 1883
rect 26 1815 108 1849
rect 26 1781 50 1815
rect 84 1781 108 1815
rect 26 1747 108 1781
rect 26 1713 50 1747
rect 84 1713 108 1747
rect 26 1679 108 1713
rect 26 1645 50 1679
rect 84 1645 108 1679
rect 26 1611 108 1645
rect 26 1577 50 1611
rect 84 1577 108 1611
rect 26 1543 108 1577
rect 26 1509 50 1543
rect 84 1509 108 1543
rect 26 1475 108 1509
rect 26 1441 50 1475
rect 84 1441 108 1475
rect 26 1407 108 1441
rect 26 1373 50 1407
rect 84 1373 108 1407
rect 26 1339 108 1373
rect 26 1305 50 1339
rect 84 1305 108 1339
rect 26 1271 108 1305
rect 26 1237 50 1271
rect 84 1237 108 1271
rect 26 1203 108 1237
rect 26 1169 50 1203
rect 84 1169 108 1203
rect 26 1135 108 1169
rect 26 1101 50 1135
rect 84 1101 108 1135
rect 26 1067 108 1101
rect 26 1033 50 1067
rect 84 1033 108 1067
rect 26 999 108 1033
rect 26 965 50 999
rect 84 965 108 999
rect 26 931 108 965
rect 26 897 50 931
rect 84 897 108 931
rect 26 863 108 897
rect 26 829 50 863
rect 84 829 108 863
rect 26 795 108 829
rect 26 761 50 795
rect 84 761 108 795
rect 26 727 108 761
rect 26 693 50 727
rect 84 693 108 727
rect 26 659 108 693
rect 26 625 50 659
rect 84 625 108 659
rect 26 591 108 625
rect 26 557 50 591
rect 84 557 108 591
rect 26 523 108 557
rect 26 489 50 523
rect 84 489 108 523
rect 26 455 108 489
rect 26 421 50 455
rect 84 421 108 455
rect 26 387 108 421
rect 26 353 50 387
rect 84 353 108 387
rect 26 319 108 353
rect 26 285 50 319
rect 84 285 108 319
rect 26 251 108 285
rect 654 2714 1538 2738
rect 654 2680 678 2714
rect 712 2680 773 2714
rect 807 2680 841 2714
rect 875 2680 909 2714
rect 943 2680 977 2714
rect 1011 2680 1045 2714
rect 1079 2680 1113 2714
rect 1147 2680 1181 2714
rect 1215 2680 1249 2714
rect 1283 2680 1317 2714
rect 1351 2680 1385 2714
rect 1419 2680 1480 2714
rect 1514 2680 1538 2714
rect 654 2656 1538 2680
rect 654 2631 736 2656
rect 654 2597 678 2631
rect 712 2597 736 2631
rect 654 2563 736 2597
rect 654 2529 678 2563
rect 712 2529 736 2563
rect 654 2495 736 2529
rect 1456 2631 1538 2656
rect 1456 2597 1480 2631
rect 1514 2597 1538 2631
rect 1456 2563 1538 2597
rect 1456 2529 1480 2563
rect 1514 2529 1538 2563
rect 654 2461 678 2495
rect 712 2461 736 2495
rect 654 2427 736 2461
rect 654 2393 678 2427
rect 712 2393 736 2427
rect 654 2359 736 2393
rect 654 2325 678 2359
rect 712 2325 736 2359
rect 654 2291 736 2325
rect 654 2257 678 2291
rect 712 2257 736 2291
rect 654 2223 736 2257
rect 654 2189 678 2223
rect 712 2189 736 2223
rect 654 2155 736 2189
rect 654 2121 678 2155
rect 712 2121 736 2155
rect 654 2087 736 2121
rect 654 2053 678 2087
rect 712 2053 736 2087
rect 654 2019 736 2053
rect 654 1985 678 2019
rect 712 1985 736 2019
rect 654 1951 736 1985
rect 654 1917 678 1951
rect 712 1917 736 1951
rect 654 1883 736 1917
rect 654 1849 678 1883
rect 712 1849 736 1883
rect 654 1815 736 1849
rect 654 1781 678 1815
rect 712 1781 736 1815
rect 654 1747 736 1781
rect 654 1713 678 1747
rect 712 1713 736 1747
rect 654 1679 736 1713
rect 654 1645 678 1679
rect 712 1645 736 1679
rect 654 1611 736 1645
rect 654 1577 678 1611
rect 712 1577 736 1611
rect 654 1543 736 1577
rect 654 1509 678 1543
rect 712 1509 736 1543
rect 654 1475 736 1509
rect 654 1441 678 1475
rect 712 1441 736 1475
rect 654 1407 736 1441
rect 654 1373 678 1407
rect 712 1373 736 1407
rect 654 1339 736 1373
rect 654 1305 678 1339
rect 712 1305 736 1339
rect 654 1271 736 1305
rect 654 1237 678 1271
rect 712 1237 736 1271
rect 654 1203 736 1237
rect 654 1169 678 1203
rect 712 1169 736 1203
rect 654 1135 736 1169
rect 654 1101 678 1135
rect 712 1101 736 1135
rect 654 1067 736 1101
rect 654 1033 678 1067
rect 712 1033 736 1067
rect 654 999 736 1033
rect 654 965 678 999
rect 712 965 736 999
rect 654 931 736 965
rect 654 897 678 931
rect 712 897 736 931
rect 654 863 736 897
rect 1456 2495 1538 2529
rect 1456 2461 1480 2495
rect 1514 2461 1538 2495
rect 1456 2427 1538 2461
rect 1456 2393 1480 2427
rect 1514 2393 1538 2427
rect 1456 2359 1538 2393
rect 1456 2325 1480 2359
rect 1514 2325 1538 2359
rect 1456 2291 1538 2325
rect 1456 2257 1480 2291
rect 1514 2257 1538 2291
rect 1456 2223 1538 2257
rect 1456 2189 1480 2223
rect 1514 2189 1538 2223
rect 1456 2155 1538 2189
rect 1456 2121 1480 2155
rect 1514 2121 1538 2155
rect 1456 2087 1538 2121
rect 1456 2053 1480 2087
rect 1514 2053 1538 2087
rect 1456 2019 1538 2053
rect 1456 1985 1480 2019
rect 1514 1985 1538 2019
rect 1456 1951 1538 1985
rect 1456 1917 1480 1951
rect 1514 1917 1538 1951
rect 1456 1883 1538 1917
rect 1456 1849 1480 1883
rect 1514 1849 1538 1883
rect 1456 1815 1538 1849
rect 1456 1781 1480 1815
rect 1514 1781 1538 1815
rect 1456 1747 1538 1781
rect 1456 1713 1480 1747
rect 1514 1713 1538 1747
rect 1456 1679 1538 1713
rect 1456 1645 1480 1679
rect 1514 1645 1538 1679
rect 1456 1611 1538 1645
rect 1456 1577 1480 1611
rect 1514 1577 1538 1611
rect 1456 1543 1538 1577
rect 1456 1509 1480 1543
rect 1514 1509 1538 1543
rect 1456 1475 1538 1509
rect 1456 1441 1480 1475
rect 1514 1441 1538 1475
rect 1456 1407 1538 1441
rect 1456 1373 1480 1407
rect 1514 1373 1538 1407
rect 1456 1339 1538 1373
rect 1456 1305 1480 1339
rect 1514 1305 1538 1339
rect 1456 1271 1538 1305
rect 1456 1237 1480 1271
rect 1514 1237 1538 1271
rect 1456 1203 1538 1237
rect 1456 1169 1480 1203
rect 1514 1169 1538 1203
rect 1456 1135 1538 1169
rect 1456 1101 1480 1135
rect 1514 1101 1538 1135
rect 1456 1067 1538 1101
rect 1456 1033 1480 1067
rect 1514 1033 1538 1067
rect 1456 999 1538 1033
rect 1456 965 1480 999
rect 1514 965 1538 999
rect 1456 931 1538 965
rect 1456 897 1480 931
rect 1514 897 1538 931
rect 654 829 678 863
rect 712 829 736 863
rect 654 795 736 829
rect 654 761 678 795
rect 712 761 736 795
rect 654 736 736 761
rect 1456 863 1538 897
rect 1456 829 1480 863
rect 1514 829 1538 863
rect 1456 795 1538 829
rect 1456 761 1480 795
rect 1514 761 1538 795
rect 1456 736 1538 761
rect 654 712 1538 736
rect 654 678 678 712
rect 712 678 773 712
rect 807 678 841 712
rect 875 678 909 712
rect 943 678 977 712
rect 1011 678 1045 712
rect 1079 678 1113 712
rect 1147 678 1181 712
rect 1215 678 1249 712
rect 1283 678 1317 712
rect 1351 678 1385 712
rect 1419 678 1480 712
rect 1514 678 1538 712
rect 654 654 1538 678
rect 2084 3107 2166 3141
rect 2084 3073 2108 3107
rect 2142 3073 2166 3107
rect 2084 3039 2166 3073
rect 2084 3005 2108 3039
rect 2142 3005 2166 3039
rect 2084 2971 2166 3005
rect 2084 2937 2108 2971
rect 2142 2937 2166 2971
rect 2084 2903 2166 2937
rect 2084 2869 2108 2903
rect 2142 2869 2166 2903
rect 2084 2835 2166 2869
rect 2084 2801 2108 2835
rect 2142 2801 2166 2835
rect 2084 2767 2166 2801
rect 2084 2733 2108 2767
rect 2142 2733 2166 2767
rect 2084 2699 2166 2733
rect 2084 2665 2108 2699
rect 2142 2665 2166 2699
rect 2084 2631 2166 2665
rect 2084 2597 2108 2631
rect 2142 2597 2166 2631
rect 2084 2563 2166 2597
rect 2084 2529 2108 2563
rect 2142 2529 2166 2563
rect 2084 2495 2166 2529
rect 2084 2461 2108 2495
rect 2142 2461 2166 2495
rect 2084 2427 2166 2461
rect 2084 2393 2108 2427
rect 2142 2393 2166 2427
rect 2084 2359 2166 2393
rect 2084 2325 2108 2359
rect 2142 2325 2166 2359
rect 2084 2291 2166 2325
rect 2084 2257 2108 2291
rect 2142 2257 2166 2291
rect 2084 2223 2166 2257
rect 2084 2189 2108 2223
rect 2142 2189 2166 2223
rect 2084 2155 2166 2189
rect 2084 2121 2108 2155
rect 2142 2121 2166 2155
rect 2084 2087 2166 2121
rect 2084 2053 2108 2087
rect 2142 2053 2166 2087
rect 2084 2019 2166 2053
rect 2084 1985 2108 2019
rect 2142 1985 2166 2019
rect 2084 1951 2166 1985
rect 2084 1917 2108 1951
rect 2142 1917 2166 1951
rect 2084 1883 2166 1917
rect 2084 1849 2108 1883
rect 2142 1849 2166 1883
rect 2084 1815 2166 1849
rect 2084 1781 2108 1815
rect 2142 1781 2166 1815
rect 2084 1747 2166 1781
rect 2084 1713 2108 1747
rect 2142 1713 2166 1747
rect 2084 1679 2166 1713
rect 2084 1645 2108 1679
rect 2142 1645 2166 1679
rect 2084 1611 2166 1645
rect 2084 1577 2108 1611
rect 2142 1577 2166 1611
rect 2084 1543 2166 1577
rect 2084 1509 2108 1543
rect 2142 1509 2166 1543
rect 2084 1475 2166 1509
rect 2084 1441 2108 1475
rect 2142 1441 2166 1475
rect 2084 1407 2166 1441
rect 2084 1373 2108 1407
rect 2142 1373 2166 1407
rect 2084 1339 2166 1373
rect 2084 1305 2108 1339
rect 2142 1305 2166 1339
rect 2084 1271 2166 1305
rect 2084 1237 2108 1271
rect 2142 1237 2166 1271
rect 2084 1203 2166 1237
rect 2084 1169 2108 1203
rect 2142 1169 2166 1203
rect 2084 1135 2166 1169
rect 2084 1101 2108 1135
rect 2142 1101 2166 1135
rect 2084 1067 2166 1101
rect 2084 1033 2108 1067
rect 2142 1033 2166 1067
rect 2084 999 2166 1033
rect 2084 965 2108 999
rect 2142 965 2166 999
rect 2084 931 2166 965
rect 2084 897 2108 931
rect 2142 897 2166 931
rect 2084 863 2166 897
rect 2084 829 2108 863
rect 2142 829 2166 863
rect 2084 795 2166 829
rect 2084 761 2108 795
rect 2142 761 2166 795
rect 2084 727 2166 761
rect 2084 693 2108 727
rect 2142 693 2166 727
rect 2084 659 2166 693
rect 2084 625 2108 659
rect 2142 625 2166 659
rect 2084 591 2166 625
rect 2084 557 2108 591
rect 2142 557 2166 591
rect 2084 523 2166 557
rect 2084 489 2108 523
rect 2142 489 2166 523
rect 2084 455 2166 489
rect 2084 421 2108 455
rect 2142 421 2166 455
rect 2084 387 2166 421
rect 2084 353 2108 387
rect 2142 353 2166 387
rect 2084 319 2166 353
rect 2084 285 2108 319
rect 2142 285 2166 319
rect 26 217 50 251
rect 84 217 108 251
rect 26 183 108 217
rect 26 149 50 183
rect 84 149 108 183
rect 26 108 108 149
rect 2084 251 2166 285
rect 2084 217 2108 251
rect 2142 217 2166 251
rect 2084 183 2166 217
rect 2084 149 2108 183
rect 2142 149 2166 183
rect 2084 108 2166 149
rect 26 84 2166 108
rect 26 50 50 84
rect 84 50 127 84
rect 161 50 195 84
rect 229 50 263 84
rect 297 50 331 84
rect 365 50 399 84
rect 433 50 467 84
rect 501 50 535 84
rect 569 50 603 84
rect 637 50 671 84
rect 705 50 739 84
rect 773 50 807 84
rect 841 50 875 84
rect 909 50 943 84
rect 977 50 1011 84
rect 1045 50 1079 84
rect 1113 50 1147 84
rect 1181 50 1215 84
rect 1249 50 1283 84
rect 1317 50 1351 84
rect 1385 50 1419 84
rect 1453 50 1487 84
rect 1521 50 1555 84
rect 1589 50 1623 84
rect 1657 50 1691 84
rect 1725 50 1759 84
rect 1793 50 1827 84
rect 1861 50 1895 84
rect 1929 50 1963 84
rect 1997 50 2031 84
rect 2065 50 2108 84
rect 2142 50 2166 84
rect 26 26 2166 50
<< nsubdiff >>
rect 252 3116 1940 3140
rect 252 3082 276 3116
rect 310 3082 365 3116
rect 399 3082 433 3116
rect 467 3082 501 3116
rect 535 3082 569 3116
rect 603 3082 637 3116
rect 671 3082 705 3116
rect 739 3082 773 3116
rect 807 3082 841 3116
rect 875 3082 909 3116
rect 943 3082 977 3116
rect 1011 3082 1045 3116
rect 1079 3082 1113 3116
rect 1147 3082 1181 3116
rect 1215 3082 1249 3116
rect 1283 3082 1317 3116
rect 1351 3082 1385 3116
rect 1419 3082 1453 3116
rect 1487 3082 1521 3116
rect 1555 3082 1589 3116
rect 1623 3082 1657 3116
rect 1691 3082 1725 3116
rect 1759 3082 1793 3116
rect 1827 3082 1882 3116
rect 1916 3082 1940 3116
rect 252 3058 1940 3082
rect 252 3039 334 3058
rect 252 3005 276 3039
rect 310 3005 334 3039
rect 252 2971 334 3005
rect 252 2937 276 2971
rect 310 2937 334 2971
rect 252 2903 334 2937
rect 252 2869 276 2903
rect 310 2869 334 2903
rect 252 2835 334 2869
rect 252 2801 276 2835
rect 310 2801 334 2835
rect 252 2767 334 2801
rect 252 2733 276 2767
rect 310 2733 334 2767
rect 1858 3039 1940 3058
rect 1858 3005 1882 3039
rect 1916 3005 1940 3039
rect 1858 2971 1940 3005
rect 1858 2937 1882 2971
rect 1916 2937 1940 2971
rect 1858 2903 1940 2937
rect 1858 2869 1882 2903
rect 1916 2869 1940 2903
rect 1858 2835 1940 2869
rect 1858 2801 1882 2835
rect 1916 2801 1940 2835
rect 1858 2767 1940 2801
rect 252 2699 334 2733
rect 252 2665 276 2699
rect 310 2665 334 2699
rect 252 2631 334 2665
rect 252 2597 276 2631
rect 310 2597 334 2631
rect 252 2563 334 2597
rect 252 2529 276 2563
rect 310 2529 334 2563
rect 252 2495 334 2529
rect 252 2461 276 2495
rect 310 2461 334 2495
rect 252 2427 334 2461
rect 252 2393 276 2427
rect 310 2393 334 2427
rect 252 2359 334 2393
rect 252 2325 276 2359
rect 310 2325 334 2359
rect 252 2291 334 2325
rect 252 2257 276 2291
rect 310 2257 334 2291
rect 252 2223 334 2257
rect 252 2189 276 2223
rect 310 2189 334 2223
rect 252 2155 334 2189
rect 252 2121 276 2155
rect 310 2121 334 2155
rect 252 2087 334 2121
rect 252 2053 276 2087
rect 310 2053 334 2087
rect 252 2019 334 2053
rect 252 1985 276 2019
rect 310 1985 334 2019
rect 252 1951 334 1985
rect 252 1917 276 1951
rect 310 1917 334 1951
rect 252 1883 334 1917
rect 252 1849 276 1883
rect 310 1849 334 1883
rect 252 1815 334 1849
rect 252 1781 276 1815
rect 310 1781 334 1815
rect 252 1747 334 1781
rect 252 1713 276 1747
rect 310 1713 334 1747
rect 252 1679 334 1713
rect 252 1645 276 1679
rect 310 1645 334 1679
rect 252 1611 334 1645
rect 252 1577 276 1611
rect 310 1577 334 1611
rect 252 1543 334 1577
rect 252 1509 276 1543
rect 310 1509 334 1543
rect 252 1475 334 1509
rect 252 1441 276 1475
rect 310 1441 334 1475
rect 252 1407 334 1441
rect 252 1373 276 1407
rect 310 1373 334 1407
rect 252 1339 334 1373
rect 252 1305 276 1339
rect 310 1305 334 1339
rect 252 1271 334 1305
rect 252 1237 276 1271
rect 310 1237 334 1271
rect 252 1203 334 1237
rect 252 1169 276 1203
rect 310 1169 334 1203
rect 252 1135 334 1169
rect 252 1101 276 1135
rect 310 1101 334 1135
rect 252 1067 334 1101
rect 252 1033 276 1067
rect 310 1033 334 1067
rect 252 999 334 1033
rect 252 965 276 999
rect 310 965 334 999
rect 252 931 334 965
rect 252 897 276 931
rect 310 897 334 931
rect 252 863 334 897
rect 252 829 276 863
rect 310 829 334 863
rect 252 795 334 829
rect 252 761 276 795
rect 310 761 334 795
rect 252 727 334 761
rect 252 693 276 727
rect 310 693 334 727
rect 252 659 334 693
rect 252 625 276 659
rect 310 625 334 659
rect 1858 2733 1882 2767
rect 1916 2733 1940 2767
rect 1858 2699 1940 2733
rect 1858 2665 1882 2699
rect 1916 2665 1940 2699
rect 1858 2631 1940 2665
rect 1858 2597 1882 2631
rect 1916 2597 1940 2631
rect 1858 2563 1940 2597
rect 1858 2529 1882 2563
rect 1916 2529 1940 2563
rect 1858 2495 1940 2529
rect 1858 2461 1882 2495
rect 1916 2461 1940 2495
rect 1858 2427 1940 2461
rect 1858 2393 1882 2427
rect 1916 2393 1940 2427
rect 1858 2359 1940 2393
rect 1858 2325 1882 2359
rect 1916 2325 1940 2359
rect 1858 2291 1940 2325
rect 1858 2257 1882 2291
rect 1916 2257 1940 2291
rect 1858 2223 1940 2257
rect 1858 2189 1882 2223
rect 1916 2189 1940 2223
rect 1858 2155 1940 2189
rect 1858 2121 1882 2155
rect 1916 2121 1940 2155
rect 1858 2087 1940 2121
rect 1858 2053 1882 2087
rect 1916 2053 1940 2087
rect 1858 2019 1940 2053
rect 1858 1985 1882 2019
rect 1916 1985 1940 2019
rect 1858 1951 1940 1985
rect 1858 1917 1882 1951
rect 1916 1917 1940 1951
rect 1858 1883 1940 1917
rect 1858 1849 1882 1883
rect 1916 1849 1940 1883
rect 1858 1815 1940 1849
rect 1858 1781 1882 1815
rect 1916 1781 1940 1815
rect 1858 1747 1940 1781
rect 1858 1713 1882 1747
rect 1916 1713 1940 1747
rect 1858 1679 1940 1713
rect 1858 1645 1882 1679
rect 1916 1645 1940 1679
rect 1858 1611 1940 1645
rect 1858 1577 1882 1611
rect 1916 1577 1940 1611
rect 1858 1543 1940 1577
rect 1858 1509 1882 1543
rect 1916 1509 1940 1543
rect 1858 1475 1940 1509
rect 1858 1441 1882 1475
rect 1916 1441 1940 1475
rect 1858 1407 1940 1441
rect 1858 1373 1882 1407
rect 1916 1373 1940 1407
rect 1858 1339 1940 1373
rect 1858 1305 1882 1339
rect 1916 1305 1940 1339
rect 1858 1271 1940 1305
rect 1858 1237 1882 1271
rect 1916 1237 1940 1271
rect 1858 1203 1940 1237
rect 1858 1169 1882 1203
rect 1916 1169 1940 1203
rect 1858 1135 1940 1169
rect 1858 1101 1882 1135
rect 1916 1101 1940 1135
rect 1858 1067 1940 1101
rect 1858 1033 1882 1067
rect 1916 1033 1940 1067
rect 1858 999 1940 1033
rect 1858 965 1882 999
rect 1916 965 1940 999
rect 1858 931 1940 965
rect 1858 897 1882 931
rect 1916 897 1940 931
rect 1858 863 1940 897
rect 1858 829 1882 863
rect 1916 829 1940 863
rect 1858 795 1940 829
rect 1858 761 1882 795
rect 1916 761 1940 795
rect 1858 727 1940 761
rect 1858 693 1882 727
rect 1916 693 1940 727
rect 1858 659 1940 693
rect 252 591 334 625
rect 252 557 276 591
rect 310 557 334 591
rect 252 523 334 557
rect 252 489 276 523
rect 310 489 334 523
rect 252 455 334 489
rect 252 421 276 455
rect 310 421 334 455
rect 252 387 334 421
rect 252 353 276 387
rect 310 353 334 387
rect 252 334 334 353
rect 1858 625 1882 659
rect 1916 625 1940 659
rect 1858 591 1940 625
rect 1858 557 1882 591
rect 1916 557 1940 591
rect 1858 523 1940 557
rect 1858 489 1882 523
rect 1916 489 1940 523
rect 1858 455 1940 489
rect 1858 421 1882 455
rect 1916 421 1940 455
rect 1858 387 1940 421
rect 1858 353 1882 387
rect 1916 353 1940 387
rect 1858 334 1940 353
rect 252 310 1940 334
rect 252 276 276 310
rect 310 276 365 310
rect 399 276 433 310
rect 467 276 501 310
rect 535 276 569 310
rect 603 276 637 310
rect 671 276 705 310
rect 739 276 773 310
rect 807 276 841 310
rect 875 276 909 310
rect 943 276 977 310
rect 1011 276 1045 310
rect 1079 276 1113 310
rect 1147 276 1181 310
rect 1215 276 1249 310
rect 1283 276 1317 310
rect 1351 276 1385 310
rect 1419 276 1453 310
rect 1487 276 1521 310
rect 1555 276 1589 310
rect 1623 276 1657 310
rect 1691 276 1725 310
rect 1759 276 1793 310
rect 1827 276 1882 310
rect 1916 276 1940 310
rect 252 252 1940 276
<< psubdiffcont >>
rect 50 3308 84 3342
rect 127 3308 161 3342
rect 195 3308 229 3342
rect 263 3308 297 3342
rect 331 3308 365 3342
rect 399 3308 433 3342
rect 467 3308 501 3342
rect 535 3308 569 3342
rect 603 3308 637 3342
rect 671 3308 705 3342
rect 739 3308 773 3342
rect 807 3308 841 3342
rect 875 3308 909 3342
rect 943 3308 977 3342
rect 1011 3308 1045 3342
rect 1079 3308 1113 3342
rect 1147 3308 1181 3342
rect 1215 3308 1249 3342
rect 1283 3308 1317 3342
rect 1351 3308 1385 3342
rect 1419 3308 1453 3342
rect 1487 3308 1521 3342
rect 1555 3308 1589 3342
rect 1623 3308 1657 3342
rect 1691 3308 1725 3342
rect 1759 3308 1793 3342
rect 1827 3308 1861 3342
rect 1895 3308 1929 3342
rect 1963 3308 1997 3342
rect 2031 3308 2065 3342
rect 2108 3308 2142 3342
rect 50 3209 84 3243
rect 50 3141 84 3175
rect 2108 3209 2142 3243
rect 2108 3141 2142 3175
rect 50 3073 84 3107
rect 50 3005 84 3039
rect 50 2937 84 2971
rect 50 2869 84 2903
rect 50 2801 84 2835
rect 50 2733 84 2767
rect 50 2665 84 2699
rect 50 2597 84 2631
rect 50 2529 84 2563
rect 50 2461 84 2495
rect 50 2393 84 2427
rect 50 2325 84 2359
rect 50 2257 84 2291
rect 50 2189 84 2223
rect 50 2121 84 2155
rect 50 2053 84 2087
rect 50 1985 84 2019
rect 50 1917 84 1951
rect 50 1849 84 1883
rect 50 1781 84 1815
rect 50 1713 84 1747
rect 50 1645 84 1679
rect 50 1577 84 1611
rect 50 1509 84 1543
rect 50 1441 84 1475
rect 50 1373 84 1407
rect 50 1305 84 1339
rect 50 1237 84 1271
rect 50 1169 84 1203
rect 50 1101 84 1135
rect 50 1033 84 1067
rect 50 965 84 999
rect 50 897 84 931
rect 50 829 84 863
rect 50 761 84 795
rect 50 693 84 727
rect 50 625 84 659
rect 50 557 84 591
rect 50 489 84 523
rect 50 421 84 455
rect 50 353 84 387
rect 50 285 84 319
rect 678 2680 712 2714
rect 773 2680 807 2714
rect 841 2680 875 2714
rect 909 2680 943 2714
rect 977 2680 1011 2714
rect 1045 2680 1079 2714
rect 1113 2680 1147 2714
rect 1181 2680 1215 2714
rect 1249 2680 1283 2714
rect 1317 2680 1351 2714
rect 1385 2680 1419 2714
rect 1480 2680 1514 2714
rect 678 2597 712 2631
rect 678 2529 712 2563
rect 1480 2597 1514 2631
rect 1480 2529 1514 2563
rect 678 2461 712 2495
rect 678 2393 712 2427
rect 678 2325 712 2359
rect 678 2257 712 2291
rect 678 2189 712 2223
rect 678 2121 712 2155
rect 678 2053 712 2087
rect 678 1985 712 2019
rect 678 1917 712 1951
rect 678 1849 712 1883
rect 678 1781 712 1815
rect 678 1713 712 1747
rect 678 1645 712 1679
rect 678 1577 712 1611
rect 678 1509 712 1543
rect 678 1441 712 1475
rect 678 1373 712 1407
rect 678 1305 712 1339
rect 678 1237 712 1271
rect 678 1169 712 1203
rect 678 1101 712 1135
rect 678 1033 712 1067
rect 678 965 712 999
rect 678 897 712 931
rect 1480 2461 1514 2495
rect 1480 2393 1514 2427
rect 1480 2325 1514 2359
rect 1480 2257 1514 2291
rect 1480 2189 1514 2223
rect 1480 2121 1514 2155
rect 1480 2053 1514 2087
rect 1480 1985 1514 2019
rect 1480 1917 1514 1951
rect 1480 1849 1514 1883
rect 1480 1781 1514 1815
rect 1480 1713 1514 1747
rect 1480 1645 1514 1679
rect 1480 1577 1514 1611
rect 1480 1509 1514 1543
rect 1480 1441 1514 1475
rect 1480 1373 1514 1407
rect 1480 1305 1514 1339
rect 1480 1237 1514 1271
rect 1480 1169 1514 1203
rect 1480 1101 1514 1135
rect 1480 1033 1514 1067
rect 1480 965 1514 999
rect 1480 897 1514 931
rect 678 829 712 863
rect 678 761 712 795
rect 1480 829 1514 863
rect 1480 761 1514 795
rect 678 678 712 712
rect 773 678 807 712
rect 841 678 875 712
rect 909 678 943 712
rect 977 678 1011 712
rect 1045 678 1079 712
rect 1113 678 1147 712
rect 1181 678 1215 712
rect 1249 678 1283 712
rect 1317 678 1351 712
rect 1385 678 1419 712
rect 1480 678 1514 712
rect 2108 3073 2142 3107
rect 2108 3005 2142 3039
rect 2108 2937 2142 2971
rect 2108 2869 2142 2903
rect 2108 2801 2142 2835
rect 2108 2733 2142 2767
rect 2108 2665 2142 2699
rect 2108 2597 2142 2631
rect 2108 2529 2142 2563
rect 2108 2461 2142 2495
rect 2108 2393 2142 2427
rect 2108 2325 2142 2359
rect 2108 2257 2142 2291
rect 2108 2189 2142 2223
rect 2108 2121 2142 2155
rect 2108 2053 2142 2087
rect 2108 1985 2142 2019
rect 2108 1917 2142 1951
rect 2108 1849 2142 1883
rect 2108 1781 2142 1815
rect 2108 1713 2142 1747
rect 2108 1645 2142 1679
rect 2108 1577 2142 1611
rect 2108 1509 2142 1543
rect 2108 1441 2142 1475
rect 2108 1373 2142 1407
rect 2108 1305 2142 1339
rect 2108 1237 2142 1271
rect 2108 1169 2142 1203
rect 2108 1101 2142 1135
rect 2108 1033 2142 1067
rect 2108 965 2142 999
rect 2108 897 2142 931
rect 2108 829 2142 863
rect 2108 761 2142 795
rect 2108 693 2142 727
rect 2108 625 2142 659
rect 2108 557 2142 591
rect 2108 489 2142 523
rect 2108 421 2142 455
rect 2108 353 2142 387
rect 2108 285 2142 319
rect 50 217 84 251
rect 50 149 84 183
rect 2108 217 2142 251
rect 2108 149 2142 183
rect 50 50 84 84
rect 127 50 161 84
rect 195 50 229 84
rect 263 50 297 84
rect 331 50 365 84
rect 399 50 433 84
rect 467 50 501 84
rect 535 50 569 84
rect 603 50 637 84
rect 671 50 705 84
rect 739 50 773 84
rect 807 50 841 84
rect 875 50 909 84
rect 943 50 977 84
rect 1011 50 1045 84
rect 1079 50 1113 84
rect 1147 50 1181 84
rect 1215 50 1249 84
rect 1283 50 1317 84
rect 1351 50 1385 84
rect 1419 50 1453 84
rect 1487 50 1521 84
rect 1555 50 1589 84
rect 1623 50 1657 84
rect 1691 50 1725 84
rect 1759 50 1793 84
rect 1827 50 1861 84
rect 1895 50 1929 84
rect 1963 50 1997 84
rect 2031 50 2065 84
rect 2108 50 2142 84
<< nsubdiffcont >>
rect 276 3082 310 3116
rect 365 3082 399 3116
rect 433 3082 467 3116
rect 501 3082 535 3116
rect 569 3082 603 3116
rect 637 3082 671 3116
rect 705 3082 739 3116
rect 773 3082 807 3116
rect 841 3082 875 3116
rect 909 3082 943 3116
rect 977 3082 1011 3116
rect 1045 3082 1079 3116
rect 1113 3082 1147 3116
rect 1181 3082 1215 3116
rect 1249 3082 1283 3116
rect 1317 3082 1351 3116
rect 1385 3082 1419 3116
rect 1453 3082 1487 3116
rect 1521 3082 1555 3116
rect 1589 3082 1623 3116
rect 1657 3082 1691 3116
rect 1725 3082 1759 3116
rect 1793 3082 1827 3116
rect 1882 3082 1916 3116
rect 276 3005 310 3039
rect 276 2937 310 2971
rect 276 2869 310 2903
rect 276 2801 310 2835
rect 276 2733 310 2767
rect 1882 3005 1916 3039
rect 1882 2937 1916 2971
rect 1882 2869 1916 2903
rect 1882 2801 1916 2835
rect 276 2665 310 2699
rect 276 2597 310 2631
rect 276 2529 310 2563
rect 276 2461 310 2495
rect 276 2393 310 2427
rect 276 2325 310 2359
rect 276 2257 310 2291
rect 276 2189 310 2223
rect 276 2121 310 2155
rect 276 2053 310 2087
rect 276 1985 310 2019
rect 276 1917 310 1951
rect 276 1849 310 1883
rect 276 1781 310 1815
rect 276 1713 310 1747
rect 276 1645 310 1679
rect 276 1577 310 1611
rect 276 1509 310 1543
rect 276 1441 310 1475
rect 276 1373 310 1407
rect 276 1305 310 1339
rect 276 1237 310 1271
rect 276 1169 310 1203
rect 276 1101 310 1135
rect 276 1033 310 1067
rect 276 965 310 999
rect 276 897 310 931
rect 276 829 310 863
rect 276 761 310 795
rect 276 693 310 727
rect 276 625 310 659
rect 1882 2733 1916 2767
rect 1882 2665 1916 2699
rect 1882 2597 1916 2631
rect 1882 2529 1916 2563
rect 1882 2461 1916 2495
rect 1882 2393 1916 2427
rect 1882 2325 1916 2359
rect 1882 2257 1916 2291
rect 1882 2189 1916 2223
rect 1882 2121 1916 2155
rect 1882 2053 1916 2087
rect 1882 1985 1916 2019
rect 1882 1917 1916 1951
rect 1882 1849 1916 1883
rect 1882 1781 1916 1815
rect 1882 1713 1916 1747
rect 1882 1645 1916 1679
rect 1882 1577 1916 1611
rect 1882 1509 1916 1543
rect 1882 1441 1916 1475
rect 1882 1373 1916 1407
rect 1882 1305 1916 1339
rect 1882 1237 1916 1271
rect 1882 1169 1916 1203
rect 1882 1101 1916 1135
rect 1882 1033 1916 1067
rect 1882 965 1916 999
rect 1882 897 1916 931
rect 1882 829 1916 863
rect 1882 761 1916 795
rect 1882 693 1916 727
rect 276 557 310 591
rect 276 489 310 523
rect 276 421 310 455
rect 276 353 310 387
rect 1882 625 1916 659
rect 1882 557 1916 591
rect 1882 489 1916 523
rect 1882 421 1916 455
rect 1882 353 1916 387
rect 276 276 310 310
rect 365 276 399 310
rect 433 276 467 310
rect 501 276 535 310
rect 569 276 603 310
rect 637 276 671 310
rect 705 276 739 310
rect 773 276 807 310
rect 841 276 875 310
rect 909 276 943 310
rect 977 276 1011 310
rect 1045 276 1079 310
rect 1113 276 1147 310
rect 1181 276 1215 310
rect 1249 276 1283 310
rect 1317 276 1351 310
rect 1385 276 1419 310
rect 1453 276 1487 310
rect 1521 276 1555 310
rect 1589 276 1623 310
rect 1657 276 1691 310
rect 1725 276 1759 310
rect 1793 276 1827 310
rect 1882 276 1916 310
<< locali >>
rect 34 3342 2158 3358
rect 34 3308 50 3342
rect 84 3308 127 3342
rect 177 3308 195 3342
rect 249 3308 263 3342
rect 321 3308 331 3342
rect 393 3308 399 3342
rect 465 3308 467 3342
rect 501 3308 503 3342
rect 569 3308 575 3342
rect 637 3308 647 3342
rect 705 3308 719 3342
rect 773 3308 791 3342
rect 841 3308 863 3342
rect 909 3308 935 3342
rect 977 3308 1007 3342
rect 1045 3308 1079 3342
rect 1113 3308 1147 3342
rect 1185 3308 1215 3342
rect 1257 3308 1283 3342
rect 1329 3308 1351 3342
rect 1401 3308 1419 3342
rect 1473 3308 1487 3342
rect 1545 3308 1555 3342
rect 1617 3308 1623 3342
rect 1689 3308 1691 3342
rect 1725 3308 1727 3342
rect 1793 3308 1799 3342
rect 1861 3308 1871 3342
rect 1929 3308 1943 3342
rect 1997 3308 2015 3342
rect 2065 3308 2108 3342
rect 2142 3308 2158 3342
rect 34 3292 2158 3308
rect 34 3261 100 3292
rect 34 3209 50 3261
rect 84 3209 100 3261
rect 34 3189 100 3209
rect 34 3141 50 3189
rect 84 3141 100 3189
rect 34 3117 100 3141
rect 2092 3261 2158 3292
rect 2092 3209 2108 3261
rect 2142 3209 2158 3261
rect 2092 3189 2158 3209
rect 2092 3141 2108 3189
rect 2142 3141 2158 3189
rect 34 3073 50 3117
rect 84 3073 100 3117
rect 34 3045 100 3073
rect 34 3005 50 3045
rect 84 3005 100 3045
rect 34 2973 100 3005
rect 34 2937 50 2973
rect 84 2937 100 2973
rect 34 2903 100 2937
rect 34 2867 50 2903
rect 84 2867 100 2903
rect 34 2835 100 2867
rect 34 2795 50 2835
rect 84 2795 100 2835
rect 34 2767 100 2795
rect 34 2723 50 2767
rect 84 2723 100 2767
rect 34 2699 100 2723
rect 34 2651 50 2699
rect 84 2651 100 2699
rect 34 2631 100 2651
rect 34 2579 50 2631
rect 84 2579 100 2631
rect 34 2563 100 2579
rect 34 2507 50 2563
rect 84 2507 100 2563
rect 34 2495 100 2507
rect 34 2435 50 2495
rect 84 2435 100 2495
rect 34 2427 100 2435
rect 34 2363 50 2427
rect 84 2363 100 2427
rect 34 2359 100 2363
rect 34 2257 50 2359
rect 84 2257 100 2359
rect 34 2253 100 2257
rect 34 2189 50 2253
rect 84 2189 100 2253
rect 34 2181 100 2189
rect 34 2121 50 2181
rect 84 2121 100 2181
rect 34 2109 100 2121
rect 34 2053 50 2109
rect 84 2053 100 2109
rect 34 2037 100 2053
rect 34 1985 50 2037
rect 84 1985 100 2037
rect 34 1965 100 1985
rect 34 1917 50 1965
rect 84 1917 100 1965
rect 34 1893 100 1917
rect 34 1849 50 1893
rect 84 1849 100 1893
rect 34 1821 100 1849
rect 34 1781 50 1821
rect 84 1781 100 1821
rect 34 1749 100 1781
rect 34 1713 50 1749
rect 84 1713 100 1749
rect 34 1679 100 1713
rect 34 1643 50 1679
rect 84 1643 100 1679
rect 34 1611 100 1643
rect 34 1571 50 1611
rect 84 1571 100 1611
rect 34 1543 100 1571
rect 34 1499 50 1543
rect 84 1499 100 1543
rect 34 1475 100 1499
rect 34 1427 50 1475
rect 84 1427 100 1475
rect 34 1407 100 1427
rect 34 1355 50 1407
rect 84 1355 100 1407
rect 34 1339 100 1355
rect 34 1283 50 1339
rect 84 1283 100 1339
rect 34 1271 100 1283
rect 34 1211 50 1271
rect 84 1211 100 1271
rect 34 1203 100 1211
rect 34 1139 50 1203
rect 84 1139 100 1203
rect 34 1135 100 1139
rect 34 1033 50 1135
rect 84 1033 100 1135
rect 34 1029 100 1033
rect 34 965 50 1029
rect 84 965 100 1029
rect 34 957 100 965
rect 34 897 50 957
rect 84 897 100 957
rect 34 885 100 897
rect 34 829 50 885
rect 84 829 100 885
rect 34 813 100 829
rect 34 761 50 813
rect 84 761 100 813
rect 34 741 100 761
rect 34 693 50 741
rect 84 693 100 741
rect 34 669 100 693
rect 34 625 50 669
rect 84 625 100 669
rect 34 597 100 625
rect 34 557 50 597
rect 84 557 100 597
rect 34 525 100 557
rect 34 489 50 525
rect 84 489 100 525
rect 34 455 100 489
rect 34 419 50 455
rect 84 419 100 455
rect 34 387 100 419
rect 34 347 50 387
rect 84 347 100 387
rect 34 319 100 347
rect 34 275 50 319
rect 84 275 100 319
rect 34 251 100 275
rect 260 3116 1932 3132
rect 260 3082 276 3116
rect 310 3082 359 3116
rect 399 3082 431 3116
rect 467 3082 501 3116
rect 537 3082 569 3116
rect 609 3082 637 3116
rect 681 3082 705 3116
rect 753 3082 773 3116
rect 825 3082 841 3116
rect 897 3082 909 3116
rect 969 3082 977 3116
rect 1041 3082 1045 3116
rect 1147 3082 1151 3116
rect 1215 3082 1223 3116
rect 1283 3082 1295 3116
rect 1351 3082 1367 3116
rect 1419 3082 1439 3116
rect 1487 3082 1511 3116
rect 1555 3082 1583 3116
rect 1623 3082 1655 3116
rect 1691 3082 1725 3116
rect 1761 3082 1793 3116
rect 1833 3082 1882 3116
rect 1916 3082 1932 3116
rect 260 3066 1932 3082
rect 260 3039 326 3066
rect 260 2975 276 3039
rect 310 2975 326 3039
rect 260 2971 326 2975
rect 260 2869 276 2971
rect 310 2869 326 2971
rect 260 2865 326 2869
rect 260 2801 276 2865
rect 310 2801 326 2865
rect 260 2793 326 2801
rect 260 2733 276 2793
rect 310 2733 326 2793
rect 260 2721 326 2733
rect 1866 3039 1932 3066
rect 1866 2975 1882 3039
rect 1916 2975 1932 3039
rect 1866 2971 1932 2975
rect 1866 2869 1882 2971
rect 1916 2869 1932 2971
rect 1866 2865 1932 2869
rect 1866 2801 1882 2865
rect 1916 2801 1932 2865
rect 1866 2793 1932 2801
rect 1866 2733 1882 2793
rect 1916 2733 1932 2793
rect 260 2665 276 2721
rect 310 2665 326 2721
rect 260 2649 326 2665
rect 260 2597 276 2649
rect 310 2597 326 2649
rect 260 2577 326 2597
rect 260 2529 276 2577
rect 310 2529 326 2577
rect 260 2505 326 2529
rect 260 2461 276 2505
rect 310 2461 326 2505
rect 260 2433 326 2461
rect 260 2393 276 2433
rect 310 2393 326 2433
rect 260 2361 326 2393
rect 260 2325 276 2361
rect 310 2325 326 2361
rect 260 2291 326 2325
rect 260 2255 276 2291
rect 310 2255 326 2291
rect 260 2223 326 2255
rect 260 2183 276 2223
rect 310 2183 326 2223
rect 260 2155 326 2183
rect 260 2111 276 2155
rect 310 2111 326 2155
rect 260 2087 326 2111
rect 260 2039 276 2087
rect 310 2039 326 2087
rect 260 2019 326 2039
rect 260 1967 276 2019
rect 310 1967 326 2019
rect 260 1951 326 1967
rect 260 1895 276 1951
rect 310 1895 326 1951
rect 260 1883 326 1895
rect 260 1823 276 1883
rect 310 1823 326 1883
rect 260 1815 326 1823
rect 260 1751 276 1815
rect 310 1751 326 1815
rect 260 1747 326 1751
rect 260 1645 276 1747
rect 310 1645 326 1747
rect 260 1641 326 1645
rect 260 1577 276 1641
rect 310 1577 326 1641
rect 260 1569 326 1577
rect 260 1509 276 1569
rect 310 1509 326 1569
rect 260 1497 326 1509
rect 260 1441 276 1497
rect 310 1441 326 1497
rect 260 1425 326 1441
rect 260 1373 276 1425
rect 310 1373 326 1425
rect 260 1353 326 1373
rect 260 1305 276 1353
rect 310 1305 326 1353
rect 260 1281 326 1305
rect 260 1237 276 1281
rect 310 1237 326 1281
rect 260 1209 326 1237
rect 260 1169 276 1209
rect 310 1169 326 1209
rect 260 1137 326 1169
rect 260 1101 276 1137
rect 310 1101 326 1137
rect 260 1067 326 1101
rect 260 1031 276 1067
rect 310 1031 326 1067
rect 260 999 326 1031
rect 260 959 276 999
rect 310 959 326 999
rect 260 931 326 959
rect 260 887 276 931
rect 310 887 326 931
rect 260 863 326 887
rect 260 815 276 863
rect 310 815 326 863
rect 260 795 326 815
rect 260 743 276 795
rect 310 743 326 795
rect 260 727 326 743
rect 260 671 276 727
rect 310 671 326 727
rect 260 659 326 671
rect 662 2714 1530 2730
rect 662 2680 678 2714
rect 712 2680 755 2714
rect 807 2680 827 2714
rect 875 2680 899 2714
rect 943 2680 971 2714
rect 1011 2680 1043 2714
rect 1079 2680 1113 2714
rect 1149 2680 1181 2714
rect 1221 2680 1249 2714
rect 1293 2680 1317 2714
rect 1365 2680 1385 2714
rect 1437 2680 1480 2714
rect 1514 2680 1530 2714
rect 662 2664 1530 2680
rect 662 2631 728 2664
rect 662 2579 678 2631
rect 712 2579 728 2631
rect 662 2563 728 2579
rect 662 2507 678 2563
rect 712 2507 728 2563
rect 662 2495 728 2507
rect 1464 2631 1530 2664
rect 1464 2579 1480 2631
rect 1514 2579 1530 2631
rect 1464 2563 1530 2579
rect 1464 2507 1480 2563
rect 1514 2507 1530 2563
rect 662 2435 678 2495
rect 712 2435 728 2495
rect 662 2427 728 2435
rect 662 2363 678 2427
rect 712 2363 728 2427
rect 662 2359 728 2363
rect 662 2257 678 2359
rect 712 2257 728 2359
rect 662 2253 728 2257
rect 662 2189 678 2253
rect 712 2189 728 2253
rect 662 2181 728 2189
rect 662 2121 678 2181
rect 712 2121 728 2181
rect 662 2109 728 2121
rect 662 2053 678 2109
rect 712 2053 728 2109
rect 662 2037 728 2053
rect 662 1985 678 2037
rect 712 1985 728 2037
rect 662 1965 728 1985
rect 662 1917 678 1965
rect 712 1917 728 1965
rect 662 1893 728 1917
rect 662 1849 678 1893
rect 712 1849 728 1893
rect 662 1821 728 1849
rect 662 1781 678 1821
rect 712 1781 728 1821
rect 662 1749 728 1781
rect 662 1713 678 1749
rect 712 1713 728 1749
rect 662 1679 728 1713
rect 662 1643 678 1679
rect 712 1643 728 1679
rect 662 1611 728 1643
rect 662 1571 678 1611
rect 712 1571 728 1611
rect 662 1543 728 1571
rect 662 1499 678 1543
rect 712 1499 728 1543
rect 662 1475 728 1499
rect 662 1427 678 1475
rect 712 1427 728 1475
rect 662 1407 728 1427
rect 662 1355 678 1407
rect 712 1355 728 1407
rect 662 1339 728 1355
rect 662 1283 678 1339
rect 712 1283 728 1339
rect 662 1271 728 1283
rect 662 1211 678 1271
rect 712 1211 728 1271
rect 662 1203 728 1211
rect 662 1139 678 1203
rect 712 1139 728 1203
rect 662 1135 728 1139
rect 662 1033 678 1135
rect 712 1033 728 1135
rect 662 1029 728 1033
rect 662 965 678 1029
rect 712 965 728 1029
rect 662 957 728 965
rect 662 897 678 957
rect 712 897 728 957
rect 662 885 728 897
rect 893 2469 1299 2499
rect 893 2461 935 2469
rect 1257 2461 1299 2469
rect 893 931 909 2461
rect 1283 931 1299 2461
rect 893 923 935 931
rect 1257 923 1299 931
rect 893 893 1299 923
rect 1464 2495 1530 2507
rect 1464 2435 1480 2495
rect 1514 2435 1530 2495
rect 1464 2427 1530 2435
rect 1464 2363 1480 2427
rect 1514 2363 1530 2427
rect 1464 2359 1530 2363
rect 1464 2257 1480 2359
rect 1514 2257 1530 2359
rect 1464 2253 1530 2257
rect 1464 2189 1480 2253
rect 1514 2189 1530 2253
rect 1464 2181 1530 2189
rect 1464 2121 1480 2181
rect 1514 2121 1530 2181
rect 1464 2109 1530 2121
rect 1464 2053 1480 2109
rect 1514 2053 1530 2109
rect 1464 2037 1530 2053
rect 1464 1985 1480 2037
rect 1514 1985 1530 2037
rect 1464 1965 1530 1985
rect 1464 1917 1480 1965
rect 1514 1917 1530 1965
rect 1464 1893 1530 1917
rect 1464 1849 1480 1893
rect 1514 1849 1530 1893
rect 1464 1821 1530 1849
rect 1464 1781 1480 1821
rect 1514 1781 1530 1821
rect 1464 1749 1530 1781
rect 1464 1713 1480 1749
rect 1514 1713 1530 1749
rect 1464 1679 1530 1713
rect 1464 1643 1480 1679
rect 1514 1643 1530 1679
rect 1464 1611 1530 1643
rect 1464 1571 1480 1611
rect 1514 1571 1530 1611
rect 1464 1543 1530 1571
rect 1464 1499 1480 1543
rect 1514 1499 1530 1543
rect 1464 1475 1530 1499
rect 1464 1427 1480 1475
rect 1514 1427 1530 1475
rect 1464 1407 1530 1427
rect 1464 1355 1480 1407
rect 1514 1355 1530 1407
rect 1464 1339 1530 1355
rect 1464 1283 1480 1339
rect 1514 1283 1530 1339
rect 1464 1271 1530 1283
rect 1464 1211 1480 1271
rect 1514 1211 1530 1271
rect 1464 1203 1530 1211
rect 1464 1139 1480 1203
rect 1514 1139 1530 1203
rect 1464 1135 1530 1139
rect 1464 1033 1480 1135
rect 1514 1033 1530 1135
rect 1464 1029 1530 1033
rect 1464 965 1480 1029
rect 1514 965 1530 1029
rect 1464 957 1530 965
rect 1464 897 1480 957
rect 1514 897 1530 957
rect 662 829 678 885
rect 712 829 728 885
rect 662 813 728 829
rect 662 761 678 813
rect 712 761 728 813
rect 662 728 728 761
rect 1464 885 1530 897
rect 1464 829 1480 885
rect 1514 829 1530 885
rect 1464 813 1530 829
rect 1464 761 1480 813
rect 1514 761 1530 813
rect 1464 728 1530 761
rect 662 712 1530 728
rect 662 678 678 712
rect 712 678 755 712
rect 807 678 827 712
rect 875 678 899 712
rect 943 678 971 712
rect 1011 678 1043 712
rect 1079 678 1113 712
rect 1149 678 1181 712
rect 1221 678 1249 712
rect 1293 678 1317 712
rect 1365 678 1385 712
rect 1437 678 1480 712
rect 1514 678 1530 712
rect 662 662 1530 678
rect 1866 2721 1932 2733
rect 1866 2665 1882 2721
rect 1916 2665 1932 2721
rect 1866 2649 1932 2665
rect 1866 2597 1882 2649
rect 1916 2597 1932 2649
rect 1866 2577 1932 2597
rect 1866 2529 1882 2577
rect 1916 2529 1932 2577
rect 1866 2505 1932 2529
rect 1866 2461 1882 2505
rect 1916 2461 1932 2505
rect 1866 2433 1932 2461
rect 1866 2393 1882 2433
rect 1916 2393 1932 2433
rect 1866 2361 1932 2393
rect 1866 2325 1882 2361
rect 1916 2325 1932 2361
rect 1866 2291 1932 2325
rect 1866 2255 1882 2291
rect 1916 2255 1932 2291
rect 1866 2223 1932 2255
rect 1866 2183 1882 2223
rect 1916 2183 1932 2223
rect 1866 2155 1932 2183
rect 1866 2111 1882 2155
rect 1916 2111 1932 2155
rect 1866 2087 1932 2111
rect 1866 2039 1882 2087
rect 1916 2039 1932 2087
rect 1866 2019 1932 2039
rect 1866 1967 1882 2019
rect 1916 1967 1932 2019
rect 1866 1951 1932 1967
rect 1866 1895 1882 1951
rect 1916 1895 1932 1951
rect 1866 1883 1932 1895
rect 1866 1823 1882 1883
rect 1916 1823 1932 1883
rect 1866 1815 1932 1823
rect 1866 1751 1882 1815
rect 1916 1751 1932 1815
rect 1866 1747 1932 1751
rect 1866 1645 1882 1747
rect 1916 1645 1932 1747
rect 1866 1641 1932 1645
rect 1866 1577 1882 1641
rect 1916 1577 1932 1641
rect 1866 1569 1932 1577
rect 1866 1509 1882 1569
rect 1916 1509 1932 1569
rect 1866 1497 1932 1509
rect 1866 1441 1882 1497
rect 1916 1441 1932 1497
rect 1866 1425 1932 1441
rect 1866 1373 1882 1425
rect 1916 1373 1932 1425
rect 1866 1353 1932 1373
rect 1866 1305 1882 1353
rect 1916 1305 1932 1353
rect 1866 1281 1932 1305
rect 1866 1237 1882 1281
rect 1916 1237 1932 1281
rect 1866 1209 1932 1237
rect 1866 1169 1882 1209
rect 1916 1169 1932 1209
rect 1866 1137 1932 1169
rect 1866 1101 1882 1137
rect 1916 1101 1932 1137
rect 1866 1067 1932 1101
rect 1866 1031 1882 1067
rect 1916 1031 1932 1067
rect 1866 999 1932 1031
rect 1866 959 1882 999
rect 1916 959 1932 999
rect 1866 931 1932 959
rect 1866 887 1882 931
rect 1916 887 1932 931
rect 1866 863 1932 887
rect 1866 815 1882 863
rect 1916 815 1932 863
rect 1866 795 1932 815
rect 1866 743 1882 795
rect 1916 743 1932 795
rect 1866 727 1932 743
rect 1866 671 1882 727
rect 1916 671 1932 727
rect 260 599 276 659
rect 310 599 326 659
rect 260 591 326 599
rect 260 527 276 591
rect 310 527 326 591
rect 260 523 326 527
rect 260 421 276 523
rect 310 421 326 523
rect 260 417 326 421
rect 260 353 276 417
rect 310 353 326 417
rect 260 326 326 353
rect 1866 659 1932 671
rect 1866 599 1882 659
rect 1916 599 1932 659
rect 1866 591 1932 599
rect 1866 527 1882 591
rect 1916 527 1932 591
rect 1866 523 1932 527
rect 1866 421 1882 523
rect 1916 421 1932 523
rect 1866 417 1932 421
rect 1866 353 1882 417
rect 1916 353 1932 417
rect 1866 326 1932 353
rect 260 310 1932 326
rect 260 276 276 310
rect 310 276 359 310
rect 399 276 431 310
rect 467 276 501 310
rect 537 276 569 310
rect 609 276 637 310
rect 681 276 705 310
rect 753 276 773 310
rect 825 276 841 310
rect 897 276 909 310
rect 969 276 977 310
rect 1041 276 1045 310
rect 1147 276 1151 310
rect 1215 276 1223 310
rect 1283 276 1295 310
rect 1351 276 1367 310
rect 1419 276 1439 310
rect 1487 276 1511 310
rect 1555 276 1583 310
rect 1623 276 1655 310
rect 1691 276 1725 310
rect 1761 276 1793 310
rect 1833 276 1882 310
rect 1916 276 1932 310
rect 260 260 1932 276
rect 2092 3117 2158 3141
rect 2092 3073 2108 3117
rect 2142 3073 2158 3117
rect 2092 3045 2158 3073
rect 2092 3005 2108 3045
rect 2142 3005 2158 3045
rect 2092 2973 2158 3005
rect 2092 2937 2108 2973
rect 2142 2937 2158 2973
rect 2092 2903 2158 2937
rect 2092 2867 2108 2903
rect 2142 2867 2158 2903
rect 2092 2835 2158 2867
rect 2092 2795 2108 2835
rect 2142 2795 2158 2835
rect 2092 2767 2158 2795
rect 2092 2723 2108 2767
rect 2142 2723 2158 2767
rect 2092 2699 2158 2723
rect 2092 2651 2108 2699
rect 2142 2651 2158 2699
rect 2092 2631 2158 2651
rect 2092 2579 2108 2631
rect 2142 2579 2158 2631
rect 2092 2563 2158 2579
rect 2092 2507 2108 2563
rect 2142 2507 2158 2563
rect 2092 2495 2158 2507
rect 2092 2435 2108 2495
rect 2142 2435 2158 2495
rect 2092 2427 2158 2435
rect 2092 2363 2108 2427
rect 2142 2363 2158 2427
rect 2092 2359 2158 2363
rect 2092 2257 2108 2359
rect 2142 2257 2158 2359
rect 2092 2253 2158 2257
rect 2092 2189 2108 2253
rect 2142 2189 2158 2253
rect 2092 2181 2158 2189
rect 2092 2121 2108 2181
rect 2142 2121 2158 2181
rect 2092 2109 2158 2121
rect 2092 2053 2108 2109
rect 2142 2053 2158 2109
rect 2092 2037 2158 2053
rect 2092 1985 2108 2037
rect 2142 1985 2158 2037
rect 2092 1965 2158 1985
rect 2092 1917 2108 1965
rect 2142 1917 2158 1965
rect 2092 1893 2158 1917
rect 2092 1849 2108 1893
rect 2142 1849 2158 1893
rect 2092 1821 2158 1849
rect 2092 1781 2108 1821
rect 2142 1781 2158 1821
rect 2092 1749 2158 1781
rect 2092 1713 2108 1749
rect 2142 1713 2158 1749
rect 2092 1679 2158 1713
rect 2092 1643 2108 1679
rect 2142 1643 2158 1679
rect 2092 1611 2158 1643
rect 2092 1571 2108 1611
rect 2142 1571 2158 1611
rect 2092 1543 2158 1571
rect 2092 1499 2108 1543
rect 2142 1499 2158 1543
rect 2092 1475 2158 1499
rect 2092 1427 2108 1475
rect 2142 1427 2158 1475
rect 2092 1407 2158 1427
rect 2092 1355 2108 1407
rect 2142 1355 2158 1407
rect 2092 1339 2158 1355
rect 2092 1283 2108 1339
rect 2142 1283 2158 1339
rect 2092 1271 2158 1283
rect 2092 1211 2108 1271
rect 2142 1211 2158 1271
rect 2092 1203 2158 1211
rect 2092 1139 2108 1203
rect 2142 1139 2158 1203
rect 2092 1135 2158 1139
rect 2092 1033 2108 1135
rect 2142 1033 2158 1135
rect 2092 1029 2158 1033
rect 2092 965 2108 1029
rect 2142 965 2158 1029
rect 2092 957 2158 965
rect 2092 897 2108 957
rect 2142 897 2158 957
rect 2092 885 2158 897
rect 2092 829 2108 885
rect 2142 829 2158 885
rect 2092 813 2158 829
rect 2092 761 2108 813
rect 2142 761 2158 813
rect 2092 741 2158 761
rect 2092 693 2108 741
rect 2142 693 2158 741
rect 2092 669 2158 693
rect 2092 625 2108 669
rect 2142 625 2158 669
rect 2092 597 2158 625
rect 2092 557 2108 597
rect 2142 557 2158 597
rect 2092 525 2158 557
rect 2092 489 2108 525
rect 2142 489 2158 525
rect 2092 455 2158 489
rect 2092 419 2108 455
rect 2142 419 2158 455
rect 2092 387 2158 419
rect 2092 347 2108 387
rect 2142 347 2158 387
rect 2092 319 2158 347
rect 2092 275 2108 319
rect 2142 275 2158 319
rect 34 203 50 251
rect 84 203 100 251
rect 34 183 100 203
rect 34 131 50 183
rect 84 131 100 183
rect 34 100 100 131
rect 2092 251 2158 275
rect 2092 203 2108 251
rect 2142 203 2158 251
rect 2092 183 2158 203
rect 2092 131 2108 183
rect 2142 131 2158 183
rect 2092 100 2158 131
rect 34 84 2158 100
rect 34 50 50 84
rect 84 50 127 84
rect 177 50 195 84
rect 249 50 263 84
rect 321 50 331 84
rect 393 50 399 84
rect 465 50 467 84
rect 501 50 503 84
rect 569 50 575 84
rect 637 50 647 84
rect 705 50 719 84
rect 773 50 791 84
rect 841 50 863 84
rect 909 50 935 84
rect 977 50 1007 84
rect 1045 50 1079 84
rect 1113 50 1147 84
rect 1185 50 1215 84
rect 1257 50 1283 84
rect 1329 50 1351 84
rect 1401 50 1419 84
rect 1473 50 1487 84
rect 1545 50 1555 84
rect 1617 50 1623 84
rect 1689 50 1691 84
rect 1725 50 1727 84
rect 1793 50 1799 84
rect 1861 50 1871 84
rect 1929 50 1943 84
rect 1997 50 2015 84
rect 2065 50 2108 84
rect 2142 50 2158 84
rect 34 34 2158 50
<< viali >>
rect 50 3308 84 3342
rect 143 3308 161 3342
rect 161 3308 177 3342
rect 215 3308 229 3342
rect 229 3308 249 3342
rect 287 3308 297 3342
rect 297 3308 321 3342
rect 359 3308 365 3342
rect 365 3308 393 3342
rect 431 3308 433 3342
rect 433 3308 465 3342
rect 503 3308 535 3342
rect 535 3308 537 3342
rect 575 3308 603 3342
rect 603 3308 609 3342
rect 647 3308 671 3342
rect 671 3308 681 3342
rect 719 3308 739 3342
rect 739 3308 753 3342
rect 791 3308 807 3342
rect 807 3308 825 3342
rect 863 3308 875 3342
rect 875 3308 897 3342
rect 935 3308 943 3342
rect 943 3308 969 3342
rect 1007 3308 1011 3342
rect 1011 3308 1041 3342
rect 1079 3308 1113 3342
rect 1151 3308 1181 3342
rect 1181 3308 1185 3342
rect 1223 3308 1249 3342
rect 1249 3308 1257 3342
rect 1295 3308 1317 3342
rect 1317 3308 1329 3342
rect 1367 3308 1385 3342
rect 1385 3308 1401 3342
rect 1439 3308 1453 3342
rect 1453 3308 1473 3342
rect 1511 3308 1521 3342
rect 1521 3308 1545 3342
rect 1583 3308 1589 3342
rect 1589 3308 1617 3342
rect 1655 3308 1657 3342
rect 1657 3308 1689 3342
rect 1727 3308 1759 3342
rect 1759 3308 1761 3342
rect 1799 3308 1827 3342
rect 1827 3308 1833 3342
rect 1871 3308 1895 3342
rect 1895 3308 1905 3342
rect 1943 3308 1963 3342
rect 1963 3308 1977 3342
rect 2015 3308 2031 3342
rect 2031 3308 2049 3342
rect 2108 3308 2142 3342
rect 50 3243 84 3261
rect 50 3227 84 3243
rect 50 3175 84 3189
rect 50 3155 84 3175
rect 2108 3243 2142 3261
rect 2108 3227 2142 3243
rect 2108 3175 2142 3189
rect 2108 3155 2142 3175
rect 50 3107 84 3117
rect 50 3083 84 3107
rect 50 3039 84 3045
rect 50 3011 84 3039
rect 50 2971 84 2973
rect 50 2939 84 2971
rect 50 2869 84 2901
rect 50 2867 84 2869
rect 50 2801 84 2829
rect 50 2795 84 2801
rect 50 2733 84 2757
rect 50 2723 84 2733
rect 50 2665 84 2685
rect 50 2651 84 2665
rect 50 2597 84 2613
rect 50 2579 84 2597
rect 50 2529 84 2541
rect 50 2507 84 2529
rect 50 2461 84 2469
rect 50 2435 84 2461
rect 50 2393 84 2397
rect 50 2363 84 2393
rect 50 2291 84 2325
rect 50 2223 84 2253
rect 50 2219 84 2223
rect 50 2155 84 2181
rect 50 2147 84 2155
rect 50 2087 84 2109
rect 50 2075 84 2087
rect 50 2019 84 2037
rect 50 2003 84 2019
rect 50 1951 84 1965
rect 50 1931 84 1951
rect 50 1883 84 1893
rect 50 1859 84 1883
rect 50 1815 84 1821
rect 50 1787 84 1815
rect 50 1747 84 1749
rect 50 1715 84 1747
rect 50 1645 84 1677
rect 50 1643 84 1645
rect 50 1577 84 1605
rect 50 1571 84 1577
rect 50 1509 84 1533
rect 50 1499 84 1509
rect 50 1441 84 1461
rect 50 1427 84 1441
rect 50 1373 84 1389
rect 50 1355 84 1373
rect 50 1305 84 1317
rect 50 1283 84 1305
rect 50 1237 84 1245
rect 50 1211 84 1237
rect 50 1169 84 1173
rect 50 1139 84 1169
rect 50 1067 84 1101
rect 50 999 84 1029
rect 50 995 84 999
rect 50 931 84 957
rect 50 923 84 931
rect 50 863 84 885
rect 50 851 84 863
rect 50 795 84 813
rect 50 779 84 795
rect 50 727 84 741
rect 50 707 84 727
rect 50 659 84 669
rect 50 635 84 659
rect 50 591 84 597
rect 50 563 84 591
rect 50 523 84 525
rect 50 491 84 523
rect 50 421 84 453
rect 50 419 84 421
rect 50 353 84 381
rect 50 347 84 353
rect 50 285 84 309
rect 50 275 84 285
rect 276 3082 310 3116
rect 359 3082 365 3116
rect 365 3082 393 3116
rect 431 3082 433 3116
rect 433 3082 465 3116
rect 503 3082 535 3116
rect 535 3082 537 3116
rect 575 3082 603 3116
rect 603 3082 609 3116
rect 647 3082 671 3116
rect 671 3082 681 3116
rect 719 3082 739 3116
rect 739 3082 753 3116
rect 791 3082 807 3116
rect 807 3082 825 3116
rect 863 3082 875 3116
rect 875 3082 897 3116
rect 935 3082 943 3116
rect 943 3082 969 3116
rect 1007 3082 1011 3116
rect 1011 3082 1041 3116
rect 1079 3082 1113 3116
rect 1151 3082 1181 3116
rect 1181 3082 1185 3116
rect 1223 3082 1249 3116
rect 1249 3082 1257 3116
rect 1295 3082 1317 3116
rect 1317 3082 1329 3116
rect 1367 3082 1385 3116
rect 1385 3082 1401 3116
rect 1439 3082 1453 3116
rect 1453 3082 1473 3116
rect 1511 3082 1521 3116
rect 1521 3082 1545 3116
rect 1583 3082 1589 3116
rect 1589 3082 1617 3116
rect 1655 3082 1657 3116
rect 1657 3082 1689 3116
rect 1727 3082 1759 3116
rect 1759 3082 1761 3116
rect 1799 3082 1827 3116
rect 1827 3082 1833 3116
rect 1882 3082 1916 3116
rect 276 3005 310 3009
rect 276 2975 310 3005
rect 276 2903 310 2937
rect 276 2835 310 2865
rect 276 2831 310 2835
rect 276 2767 310 2793
rect 276 2759 310 2767
rect 1882 3005 1916 3009
rect 1882 2975 1916 3005
rect 1882 2903 1916 2937
rect 1882 2835 1916 2865
rect 1882 2831 1916 2835
rect 1882 2767 1916 2793
rect 1882 2759 1916 2767
rect 276 2699 310 2721
rect 276 2687 310 2699
rect 276 2631 310 2649
rect 276 2615 310 2631
rect 276 2563 310 2577
rect 276 2543 310 2563
rect 276 2495 310 2505
rect 276 2471 310 2495
rect 276 2427 310 2433
rect 276 2399 310 2427
rect 276 2359 310 2361
rect 276 2327 310 2359
rect 276 2257 310 2289
rect 276 2255 310 2257
rect 276 2189 310 2217
rect 276 2183 310 2189
rect 276 2121 310 2145
rect 276 2111 310 2121
rect 276 2053 310 2073
rect 276 2039 310 2053
rect 276 1985 310 2001
rect 276 1967 310 1985
rect 276 1917 310 1929
rect 276 1895 310 1917
rect 276 1849 310 1857
rect 276 1823 310 1849
rect 276 1781 310 1785
rect 276 1751 310 1781
rect 276 1679 310 1713
rect 276 1611 310 1641
rect 276 1607 310 1611
rect 276 1543 310 1569
rect 276 1535 310 1543
rect 276 1475 310 1497
rect 276 1463 310 1475
rect 276 1407 310 1425
rect 276 1391 310 1407
rect 276 1339 310 1353
rect 276 1319 310 1339
rect 276 1271 310 1281
rect 276 1247 310 1271
rect 276 1203 310 1209
rect 276 1175 310 1203
rect 276 1135 310 1137
rect 276 1103 310 1135
rect 276 1033 310 1065
rect 276 1031 310 1033
rect 276 965 310 993
rect 276 959 310 965
rect 276 897 310 921
rect 276 887 310 897
rect 276 829 310 849
rect 276 815 310 829
rect 276 761 310 777
rect 276 743 310 761
rect 276 693 310 705
rect 276 671 310 693
rect 678 2680 712 2714
rect 755 2680 773 2714
rect 773 2680 789 2714
rect 827 2680 841 2714
rect 841 2680 861 2714
rect 899 2680 909 2714
rect 909 2680 933 2714
rect 971 2680 977 2714
rect 977 2680 1005 2714
rect 1043 2680 1045 2714
rect 1045 2680 1077 2714
rect 1115 2680 1147 2714
rect 1147 2680 1149 2714
rect 1187 2680 1215 2714
rect 1215 2680 1221 2714
rect 1259 2680 1283 2714
rect 1283 2680 1293 2714
rect 1331 2680 1351 2714
rect 1351 2680 1365 2714
rect 1403 2680 1419 2714
rect 1419 2680 1437 2714
rect 1480 2680 1514 2714
rect 678 2597 712 2613
rect 678 2579 712 2597
rect 678 2529 712 2541
rect 678 2507 712 2529
rect 1480 2597 1514 2613
rect 1480 2579 1514 2597
rect 1480 2529 1514 2541
rect 1480 2507 1514 2529
rect 678 2461 712 2469
rect 678 2435 712 2461
rect 678 2393 712 2397
rect 678 2363 712 2393
rect 678 2291 712 2325
rect 678 2223 712 2253
rect 678 2219 712 2223
rect 678 2155 712 2181
rect 678 2147 712 2155
rect 678 2087 712 2109
rect 678 2075 712 2087
rect 678 2019 712 2037
rect 678 2003 712 2019
rect 678 1951 712 1965
rect 678 1931 712 1951
rect 678 1883 712 1893
rect 678 1859 712 1883
rect 678 1815 712 1821
rect 678 1787 712 1815
rect 678 1747 712 1749
rect 678 1715 712 1747
rect 678 1645 712 1677
rect 678 1643 712 1645
rect 678 1577 712 1605
rect 678 1571 712 1577
rect 678 1509 712 1533
rect 678 1499 712 1509
rect 678 1441 712 1461
rect 678 1427 712 1441
rect 678 1373 712 1389
rect 678 1355 712 1373
rect 678 1305 712 1317
rect 678 1283 712 1305
rect 678 1237 712 1245
rect 678 1211 712 1237
rect 678 1169 712 1173
rect 678 1139 712 1169
rect 678 1067 712 1101
rect 678 999 712 1029
rect 678 995 712 999
rect 678 931 712 957
rect 678 923 712 931
rect 935 2461 1257 2469
rect 935 931 1257 2461
rect 935 923 1257 931
rect 1480 2461 1514 2469
rect 1480 2435 1514 2461
rect 1480 2393 1514 2397
rect 1480 2363 1514 2393
rect 1480 2291 1514 2325
rect 1480 2223 1514 2253
rect 1480 2219 1514 2223
rect 1480 2155 1514 2181
rect 1480 2147 1514 2155
rect 1480 2087 1514 2109
rect 1480 2075 1514 2087
rect 1480 2019 1514 2037
rect 1480 2003 1514 2019
rect 1480 1951 1514 1965
rect 1480 1931 1514 1951
rect 1480 1883 1514 1893
rect 1480 1859 1514 1883
rect 1480 1815 1514 1821
rect 1480 1787 1514 1815
rect 1480 1747 1514 1749
rect 1480 1715 1514 1747
rect 1480 1645 1514 1677
rect 1480 1643 1514 1645
rect 1480 1577 1514 1605
rect 1480 1571 1514 1577
rect 1480 1509 1514 1533
rect 1480 1499 1514 1509
rect 1480 1441 1514 1461
rect 1480 1427 1514 1441
rect 1480 1373 1514 1389
rect 1480 1355 1514 1373
rect 1480 1305 1514 1317
rect 1480 1283 1514 1305
rect 1480 1237 1514 1245
rect 1480 1211 1514 1237
rect 1480 1169 1514 1173
rect 1480 1139 1514 1169
rect 1480 1067 1514 1101
rect 1480 999 1514 1029
rect 1480 995 1514 999
rect 1480 931 1514 957
rect 1480 923 1514 931
rect 678 863 712 885
rect 678 851 712 863
rect 678 795 712 813
rect 678 779 712 795
rect 1480 863 1514 885
rect 1480 851 1514 863
rect 1480 795 1514 813
rect 1480 779 1514 795
rect 678 678 712 712
rect 755 678 773 712
rect 773 678 789 712
rect 827 678 841 712
rect 841 678 861 712
rect 899 678 909 712
rect 909 678 933 712
rect 971 678 977 712
rect 977 678 1005 712
rect 1043 678 1045 712
rect 1045 678 1077 712
rect 1115 678 1147 712
rect 1147 678 1149 712
rect 1187 678 1215 712
rect 1215 678 1221 712
rect 1259 678 1283 712
rect 1283 678 1293 712
rect 1331 678 1351 712
rect 1351 678 1365 712
rect 1403 678 1419 712
rect 1419 678 1437 712
rect 1480 678 1514 712
rect 1882 2699 1916 2721
rect 1882 2687 1916 2699
rect 1882 2631 1916 2649
rect 1882 2615 1916 2631
rect 1882 2563 1916 2577
rect 1882 2543 1916 2563
rect 1882 2495 1916 2505
rect 1882 2471 1916 2495
rect 1882 2427 1916 2433
rect 1882 2399 1916 2427
rect 1882 2359 1916 2361
rect 1882 2327 1916 2359
rect 1882 2257 1916 2289
rect 1882 2255 1916 2257
rect 1882 2189 1916 2217
rect 1882 2183 1916 2189
rect 1882 2121 1916 2145
rect 1882 2111 1916 2121
rect 1882 2053 1916 2073
rect 1882 2039 1916 2053
rect 1882 1985 1916 2001
rect 1882 1967 1916 1985
rect 1882 1917 1916 1929
rect 1882 1895 1916 1917
rect 1882 1849 1916 1857
rect 1882 1823 1916 1849
rect 1882 1781 1916 1785
rect 1882 1751 1916 1781
rect 1882 1679 1916 1713
rect 1882 1611 1916 1641
rect 1882 1607 1916 1611
rect 1882 1543 1916 1569
rect 1882 1535 1916 1543
rect 1882 1475 1916 1497
rect 1882 1463 1916 1475
rect 1882 1407 1916 1425
rect 1882 1391 1916 1407
rect 1882 1339 1916 1353
rect 1882 1319 1916 1339
rect 1882 1271 1916 1281
rect 1882 1247 1916 1271
rect 1882 1203 1916 1209
rect 1882 1175 1916 1203
rect 1882 1135 1916 1137
rect 1882 1103 1916 1135
rect 1882 1033 1916 1065
rect 1882 1031 1916 1033
rect 1882 965 1916 993
rect 1882 959 1916 965
rect 1882 897 1916 921
rect 1882 887 1916 897
rect 1882 829 1916 849
rect 1882 815 1916 829
rect 1882 761 1916 777
rect 1882 743 1916 761
rect 1882 693 1916 705
rect 1882 671 1916 693
rect 276 625 310 633
rect 276 599 310 625
rect 276 557 310 561
rect 276 527 310 557
rect 276 455 310 489
rect 276 387 310 417
rect 276 383 310 387
rect 1882 625 1916 633
rect 1882 599 1916 625
rect 1882 557 1916 561
rect 1882 527 1916 557
rect 1882 455 1916 489
rect 1882 387 1916 417
rect 1882 383 1916 387
rect 276 276 310 310
rect 359 276 365 310
rect 365 276 393 310
rect 431 276 433 310
rect 433 276 465 310
rect 503 276 535 310
rect 535 276 537 310
rect 575 276 603 310
rect 603 276 609 310
rect 647 276 671 310
rect 671 276 681 310
rect 719 276 739 310
rect 739 276 753 310
rect 791 276 807 310
rect 807 276 825 310
rect 863 276 875 310
rect 875 276 897 310
rect 935 276 943 310
rect 943 276 969 310
rect 1007 276 1011 310
rect 1011 276 1041 310
rect 1079 276 1113 310
rect 1151 276 1181 310
rect 1181 276 1185 310
rect 1223 276 1249 310
rect 1249 276 1257 310
rect 1295 276 1317 310
rect 1317 276 1329 310
rect 1367 276 1385 310
rect 1385 276 1401 310
rect 1439 276 1453 310
rect 1453 276 1473 310
rect 1511 276 1521 310
rect 1521 276 1545 310
rect 1583 276 1589 310
rect 1589 276 1617 310
rect 1655 276 1657 310
rect 1657 276 1689 310
rect 1727 276 1759 310
rect 1759 276 1761 310
rect 1799 276 1827 310
rect 1827 276 1833 310
rect 1882 276 1916 310
rect 2108 3107 2142 3117
rect 2108 3083 2142 3107
rect 2108 3039 2142 3045
rect 2108 3011 2142 3039
rect 2108 2971 2142 2973
rect 2108 2939 2142 2971
rect 2108 2869 2142 2901
rect 2108 2867 2142 2869
rect 2108 2801 2142 2829
rect 2108 2795 2142 2801
rect 2108 2733 2142 2757
rect 2108 2723 2142 2733
rect 2108 2665 2142 2685
rect 2108 2651 2142 2665
rect 2108 2597 2142 2613
rect 2108 2579 2142 2597
rect 2108 2529 2142 2541
rect 2108 2507 2142 2529
rect 2108 2461 2142 2469
rect 2108 2435 2142 2461
rect 2108 2393 2142 2397
rect 2108 2363 2142 2393
rect 2108 2291 2142 2325
rect 2108 2223 2142 2253
rect 2108 2219 2142 2223
rect 2108 2155 2142 2181
rect 2108 2147 2142 2155
rect 2108 2087 2142 2109
rect 2108 2075 2142 2087
rect 2108 2019 2142 2037
rect 2108 2003 2142 2019
rect 2108 1951 2142 1965
rect 2108 1931 2142 1951
rect 2108 1883 2142 1893
rect 2108 1859 2142 1883
rect 2108 1815 2142 1821
rect 2108 1787 2142 1815
rect 2108 1747 2142 1749
rect 2108 1715 2142 1747
rect 2108 1645 2142 1677
rect 2108 1643 2142 1645
rect 2108 1577 2142 1605
rect 2108 1571 2142 1577
rect 2108 1509 2142 1533
rect 2108 1499 2142 1509
rect 2108 1441 2142 1461
rect 2108 1427 2142 1441
rect 2108 1373 2142 1389
rect 2108 1355 2142 1373
rect 2108 1305 2142 1317
rect 2108 1283 2142 1305
rect 2108 1237 2142 1245
rect 2108 1211 2142 1237
rect 2108 1169 2142 1173
rect 2108 1139 2142 1169
rect 2108 1067 2142 1101
rect 2108 999 2142 1029
rect 2108 995 2142 999
rect 2108 931 2142 957
rect 2108 923 2142 931
rect 2108 863 2142 885
rect 2108 851 2142 863
rect 2108 795 2142 813
rect 2108 779 2142 795
rect 2108 727 2142 741
rect 2108 707 2142 727
rect 2108 659 2142 669
rect 2108 635 2142 659
rect 2108 591 2142 597
rect 2108 563 2142 591
rect 2108 523 2142 525
rect 2108 491 2142 523
rect 2108 421 2142 453
rect 2108 419 2142 421
rect 2108 353 2142 381
rect 2108 347 2142 353
rect 2108 285 2142 309
rect 2108 275 2142 285
rect 50 217 84 237
rect 50 203 84 217
rect 50 149 84 165
rect 50 131 84 149
rect 2108 217 2142 237
rect 2108 203 2142 217
rect 2108 149 2142 165
rect 2108 131 2142 149
rect 50 50 84 84
rect 143 50 161 84
rect 161 50 177 84
rect 215 50 229 84
rect 229 50 249 84
rect 287 50 297 84
rect 297 50 321 84
rect 359 50 365 84
rect 365 50 393 84
rect 431 50 433 84
rect 433 50 465 84
rect 503 50 535 84
rect 535 50 537 84
rect 575 50 603 84
rect 603 50 609 84
rect 647 50 671 84
rect 671 50 681 84
rect 719 50 739 84
rect 739 50 753 84
rect 791 50 807 84
rect 807 50 825 84
rect 863 50 875 84
rect 875 50 897 84
rect 935 50 943 84
rect 943 50 969 84
rect 1007 50 1011 84
rect 1011 50 1041 84
rect 1079 50 1113 84
rect 1151 50 1181 84
rect 1181 50 1185 84
rect 1223 50 1249 84
rect 1249 50 1257 84
rect 1295 50 1317 84
rect 1317 50 1329 84
rect 1367 50 1385 84
rect 1385 50 1401 84
rect 1439 50 1453 84
rect 1453 50 1473 84
rect 1511 50 1521 84
rect 1521 50 1545 84
rect 1583 50 1589 84
rect 1589 50 1617 84
rect 1655 50 1657 84
rect 1657 50 1689 84
rect 1727 50 1759 84
rect 1759 50 1761 84
rect 1799 50 1827 84
rect 1827 50 1833 84
rect 1871 50 1895 84
rect 1895 50 1905 84
rect 1943 50 1963 84
rect 1963 50 1977 84
rect 2015 50 2031 84
rect 2031 50 2049 84
rect 2108 50 2142 84
<< metal1 >>
rect 38 3342 2154 3354
rect 38 3308 50 3342
rect 84 3308 143 3342
rect 177 3308 215 3342
rect 249 3308 287 3342
rect 321 3308 359 3342
rect 393 3308 431 3342
rect 465 3308 503 3342
rect 537 3308 575 3342
rect 609 3308 647 3342
rect 681 3308 719 3342
rect 753 3308 791 3342
rect 825 3308 863 3342
rect 897 3308 935 3342
rect 969 3308 1007 3342
rect 1041 3308 1079 3342
rect 1113 3308 1151 3342
rect 1185 3308 1223 3342
rect 1257 3308 1295 3342
rect 1329 3308 1367 3342
rect 1401 3308 1439 3342
rect 1473 3308 1511 3342
rect 1545 3308 1583 3342
rect 1617 3308 1655 3342
rect 1689 3308 1727 3342
rect 1761 3308 1799 3342
rect 1833 3308 1871 3342
rect 1905 3308 1943 3342
rect 1977 3308 2015 3342
rect 2049 3308 2108 3342
rect 2142 3308 2154 3342
rect 38 3296 2154 3308
rect 38 3261 96 3296
rect 38 3227 50 3261
rect 84 3227 96 3261
rect 38 3189 96 3227
rect 38 3155 50 3189
rect 84 3155 96 3189
rect 38 3117 96 3155
rect 2096 3261 2154 3296
rect 2096 3227 2108 3261
rect 2142 3227 2154 3261
rect 2096 3189 2154 3227
rect 2096 3155 2108 3189
rect 2142 3155 2154 3189
rect 38 3083 50 3117
rect 84 3083 96 3117
rect 38 3045 96 3083
rect 38 3011 50 3045
rect 84 3011 96 3045
rect 38 2973 96 3011
rect 38 2939 50 2973
rect 84 2939 96 2973
rect 38 2901 96 2939
rect 38 2867 50 2901
rect 84 2867 96 2901
rect 38 2829 96 2867
rect 38 2795 50 2829
rect 84 2795 96 2829
rect 38 2757 96 2795
rect 38 2723 50 2757
rect 84 2723 96 2757
rect 38 2685 96 2723
rect 38 2651 50 2685
rect 84 2651 96 2685
rect 38 2613 96 2651
rect 38 2579 50 2613
rect 84 2579 96 2613
rect 38 2541 96 2579
rect 38 2507 50 2541
rect 84 2507 96 2541
rect 38 2469 96 2507
rect 38 2435 50 2469
rect 84 2435 96 2469
rect 38 2397 96 2435
rect 38 2363 50 2397
rect 84 2363 96 2397
rect 38 2325 96 2363
rect 38 2291 50 2325
rect 84 2291 96 2325
rect 38 2253 96 2291
rect 38 2219 50 2253
rect 84 2219 96 2253
rect 38 2181 96 2219
rect 38 2147 50 2181
rect 84 2147 96 2181
rect 38 2109 96 2147
rect 38 2075 50 2109
rect 84 2075 96 2109
rect 38 2037 96 2075
rect 38 2003 50 2037
rect 84 2003 96 2037
rect 38 1965 96 2003
rect 38 1931 50 1965
rect 84 1931 96 1965
rect 38 1893 96 1931
rect 38 1859 50 1893
rect 84 1859 96 1893
rect 38 1821 96 1859
rect 38 1787 50 1821
rect 84 1787 96 1821
rect 38 1749 96 1787
rect 38 1715 50 1749
rect 84 1715 96 1749
rect 38 1677 96 1715
rect 38 1643 50 1677
rect 84 1643 96 1677
rect 38 1605 96 1643
rect 38 1571 50 1605
rect 84 1571 96 1605
rect 38 1533 96 1571
rect 38 1499 50 1533
rect 84 1499 96 1533
rect 38 1461 96 1499
rect 38 1427 50 1461
rect 84 1427 96 1461
rect 38 1389 96 1427
rect 38 1355 50 1389
rect 84 1355 96 1389
rect 38 1317 96 1355
rect 38 1283 50 1317
rect 84 1283 96 1317
rect 38 1245 96 1283
rect 38 1211 50 1245
rect 84 1211 96 1245
rect 38 1173 96 1211
rect 38 1139 50 1173
rect 84 1139 96 1173
rect 38 1101 96 1139
rect 38 1067 50 1101
rect 84 1067 96 1101
rect 38 1029 96 1067
rect 38 995 50 1029
rect 84 995 96 1029
rect 38 957 96 995
rect 38 923 50 957
rect 84 923 96 957
rect 38 885 96 923
rect 38 851 50 885
rect 84 851 96 885
rect 38 813 96 851
rect 38 779 50 813
rect 84 779 96 813
rect 38 741 96 779
rect 38 707 50 741
rect 84 707 96 741
rect 38 669 96 707
rect 38 635 50 669
rect 84 635 96 669
rect 38 597 96 635
rect 38 563 50 597
rect 84 563 96 597
rect 38 525 96 563
rect 38 491 50 525
rect 84 491 96 525
rect 38 453 96 491
rect 38 419 50 453
rect 84 419 96 453
rect 38 381 96 419
rect 38 347 50 381
rect 84 347 96 381
rect 38 309 96 347
rect 38 275 50 309
rect 84 275 96 309
rect 38 237 96 275
rect 264 3116 1928 3128
rect 264 3082 276 3116
rect 310 3082 359 3116
rect 393 3082 431 3116
rect 465 3082 503 3116
rect 537 3082 575 3116
rect 609 3082 647 3116
rect 681 3082 719 3116
rect 753 3082 791 3116
rect 825 3082 863 3116
rect 897 3082 935 3116
rect 969 3082 1007 3116
rect 1041 3082 1079 3116
rect 1113 3082 1151 3116
rect 1185 3082 1223 3116
rect 1257 3082 1295 3116
rect 1329 3082 1367 3116
rect 1401 3082 1439 3116
rect 1473 3082 1511 3116
rect 1545 3082 1583 3116
rect 1617 3082 1655 3116
rect 1689 3082 1727 3116
rect 1761 3082 1799 3116
rect 1833 3082 1882 3116
rect 1916 3082 1928 3116
rect 264 3070 1928 3082
rect 264 3009 322 3070
rect 264 2975 276 3009
rect 310 2975 322 3009
rect 264 2937 322 2975
rect 264 2903 276 2937
rect 310 2903 322 2937
rect 264 2865 322 2903
rect 264 2831 276 2865
rect 310 2831 322 2865
rect 264 2793 322 2831
rect 264 2759 276 2793
rect 310 2759 322 2793
rect 264 2721 322 2759
rect 1870 3009 1928 3070
rect 1870 2975 1882 3009
rect 1916 2975 1928 3009
rect 1870 2937 1928 2975
rect 1870 2903 1882 2937
rect 1916 2903 1928 2937
rect 1870 2865 1928 2903
rect 1870 2831 1882 2865
rect 1916 2831 1928 2865
rect 1870 2793 1928 2831
rect 1870 2759 1882 2793
rect 1916 2759 1928 2793
rect 264 2687 276 2721
rect 310 2687 322 2721
rect 264 2649 322 2687
rect 264 2615 276 2649
rect 310 2615 322 2649
rect 264 2577 322 2615
rect 264 2543 276 2577
rect 310 2543 322 2577
rect 264 2505 322 2543
rect 264 2471 276 2505
rect 310 2471 322 2505
rect 264 2433 322 2471
rect 264 2399 276 2433
rect 310 2399 322 2433
rect 264 2361 322 2399
rect 264 2327 276 2361
rect 310 2327 322 2361
rect 264 2289 322 2327
rect 264 2255 276 2289
rect 310 2255 322 2289
rect 264 2217 322 2255
rect 264 2183 276 2217
rect 310 2183 322 2217
rect 264 2145 322 2183
rect 264 2111 276 2145
rect 310 2111 322 2145
rect 264 2073 322 2111
rect 264 2039 276 2073
rect 310 2039 322 2073
rect 264 2001 322 2039
rect 264 1967 276 2001
rect 310 1967 322 2001
rect 264 1929 322 1967
rect 264 1895 276 1929
rect 310 1895 322 1929
rect 264 1857 322 1895
rect 264 1823 276 1857
rect 310 1823 322 1857
rect 264 1785 322 1823
rect 264 1751 276 1785
rect 310 1751 322 1785
rect 264 1713 322 1751
rect 264 1679 276 1713
rect 310 1679 322 1713
rect 264 1641 322 1679
rect 264 1607 276 1641
rect 310 1607 322 1641
rect 264 1569 322 1607
rect 264 1535 276 1569
rect 310 1535 322 1569
rect 264 1497 322 1535
rect 264 1463 276 1497
rect 310 1463 322 1497
rect 264 1425 322 1463
rect 264 1391 276 1425
rect 310 1391 322 1425
rect 264 1353 322 1391
rect 264 1319 276 1353
rect 310 1319 322 1353
rect 264 1281 322 1319
rect 264 1247 276 1281
rect 310 1247 322 1281
rect 264 1209 322 1247
rect 264 1175 276 1209
rect 310 1175 322 1209
rect 264 1137 322 1175
rect 264 1103 276 1137
rect 310 1103 322 1137
rect 264 1065 322 1103
rect 264 1031 276 1065
rect 310 1031 322 1065
rect 264 993 322 1031
rect 264 959 276 993
rect 310 959 322 993
rect 264 921 322 959
rect 264 887 276 921
rect 310 887 322 921
rect 264 849 322 887
rect 264 815 276 849
rect 310 815 322 849
rect 264 777 322 815
rect 264 743 276 777
rect 310 743 322 777
rect 264 705 322 743
rect 264 671 276 705
rect 310 671 322 705
rect 264 633 322 671
rect 666 2714 1526 2726
rect 666 2680 678 2714
rect 712 2680 755 2714
rect 789 2680 827 2714
rect 861 2680 899 2714
rect 933 2680 971 2714
rect 1005 2680 1043 2714
rect 1077 2680 1115 2714
rect 1149 2680 1187 2714
rect 1221 2680 1259 2714
rect 1293 2680 1331 2714
rect 1365 2680 1403 2714
rect 1437 2680 1480 2714
rect 1514 2680 1526 2714
rect 666 2668 1526 2680
rect 666 2613 724 2668
rect 666 2579 678 2613
rect 712 2579 724 2613
rect 666 2541 724 2579
rect 666 2507 678 2541
rect 712 2507 724 2541
rect 666 2469 724 2507
rect 1468 2613 1526 2668
rect 1468 2579 1480 2613
rect 1514 2579 1526 2613
rect 1468 2541 1526 2579
rect 1468 2507 1480 2541
rect 1514 2507 1526 2541
rect 666 2435 678 2469
rect 712 2435 724 2469
rect 666 2397 724 2435
rect 666 2363 678 2397
rect 712 2363 724 2397
rect 666 2325 724 2363
rect 666 2291 678 2325
rect 712 2291 724 2325
rect 666 2253 724 2291
rect 666 2219 678 2253
rect 712 2219 724 2253
rect 666 2181 724 2219
rect 666 2147 678 2181
rect 712 2147 724 2181
rect 666 2109 724 2147
rect 666 2075 678 2109
rect 712 2075 724 2109
rect 666 2037 724 2075
rect 666 2003 678 2037
rect 712 2003 724 2037
rect 666 1965 724 2003
rect 666 1931 678 1965
rect 712 1931 724 1965
rect 666 1893 724 1931
rect 666 1859 678 1893
rect 712 1859 724 1893
rect 666 1821 724 1859
rect 666 1787 678 1821
rect 712 1787 724 1821
rect 666 1749 724 1787
rect 666 1715 678 1749
rect 712 1715 724 1749
rect 666 1677 724 1715
rect 666 1643 678 1677
rect 712 1643 724 1677
rect 666 1605 724 1643
rect 666 1571 678 1605
rect 712 1571 724 1605
rect 666 1533 724 1571
rect 666 1499 678 1533
rect 712 1499 724 1533
rect 666 1461 724 1499
rect 666 1427 678 1461
rect 712 1427 724 1461
rect 666 1389 724 1427
rect 666 1355 678 1389
rect 712 1355 724 1389
rect 666 1317 724 1355
rect 666 1283 678 1317
rect 712 1283 724 1317
rect 666 1245 724 1283
rect 666 1211 678 1245
rect 712 1211 724 1245
rect 666 1173 724 1211
rect 666 1139 678 1173
rect 712 1139 724 1173
rect 666 1101 724 1139
rect 666 1067 678 1101
rect 712 1067 724 1101
rect 666 1029 724 1067
rect 666 995 678 1029
rect 712 995 724 1029
rect 666 957 724 995
rect 666 923 678 957
rect 712 923 724 957
rect 666 885 724 923
rect 923 2469 1269 2481
rect 923 923 935 2469
rect 1257 923 1269 2469
rect 923 911 1269 923
rect 1468 2469 1526 2507
rect 1468 2435 1480 2469
rect 1514 2435 1526 2469
rect 1468 2397 1526 2435
rect 1468 2363 1480 2397
rect 1514 2363 1526 2397
rect 1468 2325 1526 2363
rect 1468 2291 1480 2325
rect 1514 2291 1526 2325
rect 1468 2253 1526 2291
rect 1468 2219 1480 2253
rect 1514 2219 1526 2253
rect 1468 2181 1526 2219
rect 1468 2147 1480 2181
rect 1514 2147 1526 2181
rect 1468 2109 1526 2147
rect 1468 2075 1480 2109
rect 1514 2075 1526 2109
rect 1468 2037 1526 2075
rect 1468 2003 1480 2037
rect 1514 2003 1526 2037
rect 1468 1965 1526 2003
rect 1468 1931 1480 1965
rect 1514 1931 1526 1965
rect 1468 1893 1526 1931
rect 1468 1859 1480 1893
rect 1514 1859 1526 1893
rect 1468 1821 1526 1859
rect 1468 1787 1480 1821
rect 1514 1787 1526 1821
rect 1468 1749 1526 1787
rect 1468 1715 1480 1749
rect 1514 1715 1526 1749
rect 1468 1677 1526 1715
rect 1468 1643 1480 1677
rect 1514 1643 1526 1677
rect 1468 1605 1526 1643
rect 1468 1571 1480 1605
rect 1514 1571 1526 1605
rect 1468 1533 1526 1571
rect 1468 1499 1480 1533
rect 1514 1499 1526 1533
rect 1468 1461 1526 1499
rect 1468 1427 1480 1461
rect 1514 1427 1526 1461
rect 1468 1389 1526 1427
rect 1468 1355 1480 1389
rect 1514 1355 1526 1389
rect 1468 1317 1526 1355
rect 1468 1283 1480 1317
rect 1514 1283 1526 1317
rect 1468 1245 1526 1283
rect 1468 1211 1480 1245
rect 1514 1211 1526 1245
rect 1468 1173 1526 1211
rect 1468 1139 1480 1173
rect 1514 1139 1526 1173
rect 1468 1101 1526 1139
rect 1468 1067 1480 1101
rect 1514 1067 1526 1101
rect 1468 1029 1526 1067
rect 1468 995 1480 1029
rect 1514 995 1526 1029
rect 1468 957 1526 995
rect 1468 923 1480 957
rect 1514 923 1526 957
rect 666 851 678 885
rect 712 851 724 885
rect 666 813 724 851
rect 666 779 678 813
rect 712 779 724 813
rect 666 724 724 779
rect 1468 885 1526 923
rect 1468 851 1480 885
rect 1514 851 1526 885
rect 1468 813 1526 851
rect 1468 779 1480 813
rect 1514 779 1526 813
rect 1468 724 1526 779
rect 666 712 1526 724
rect 666 678 678 712
rect 712 678 755 712
rect 789 678 827 712
rect 861 678 899 712
rect 933 678 971 712
rect 1005 678 1043 712
rect 1077 678 1115 712
rect 1149 678 1187 712
rect 1221 678 1259 712
rect 1293 678 1331 712
rect 1365 678 1403 712
rect 1437 678 1480 712
rect 1514 678 1526 712
rect 666 666 1526 678
rect 1870 2721 1928 2759
rect 1870 2687 1882 2721
rect 1916 2687 1928 2721
rect 1870 2649 1928 2687
rect 1870 2615 1882 2649
rect 1916 2615 1928 2649
rect 1870 2577 1928 2615
rect 1870 2543 1882 2577
rect 1916 2543 1928 2577
rect 1870 2505 1928 2543
rect 1870 2471 1882 2505
rect 1916 2471 1928 2505
rect 1870 2433 1928 2471
rect 1870 2399 1882 2433
rect 1916 2399 1928 2433
rect 1870 2361 1928 2399
rect 1870 2327 1882 2361
rect 1916 2327 1928 2361
rect 1870 2289 1928 2327
rect 1870 2255 1882 2289
rect 1916 2255 1928 2289
rect 1870 2217 1928 2255
rect 1870 2183 1882 2217
rect 1916 2183 1928 2217
rect 1870 2145 1928 2183
rect 1870 2111 1882 2145
rect 1916 2111 1928 2145
rect 1870 2073 1928 2111
rect 1870 2039 1882 2073
rect 1916 2039 1928 2073
rect 1870 2001 1928 2039
rect 1870 1967 1882 2001
rect 1916 1967 1928 2001
rect 1870 1929 1928 1967
rect 1870 1895 1882 1929
rect 1916 1895 1928 1929
rect 1870 1857 1928 1895
rect 1870 1823 1882 1857
rect 1916 1823 1928 1857
rect 1870 1785 1928 1823
rect 1870 1751 1882 1785
rect 1916 1751 1928 1785
rect 1870 1713 1928 1751
rect 1870 1679 1882 1713
rect 1916 1679 1928 1713
rect 1870 1641 1928 1679
rect 1870 1607 1882 1641
rect 1916 1607 1928 1641
rect 1870 1569 1928 1607
rect 1870 1535 1882 1569
rect 1916 1535 1928 1569
rect 1870 1497 1928 1535
rect 1870 1463 1882 1497
rect 1916 1463 1928 1497
rect 1870 1425 1928 1463
rect 1870 1391 1882 1425
rect 1916 1391 1928 1425
rect 1870 1353 1928 1391
rect 1870 1319 1882 1353
rect 1916 1319 1928 1353
rect 1870 1281 1928 1319
rect 1870 1247 1882 1281
rect 1916 1247 1928 1281
rect 1870 1209 1928 1247
rect 1870 1175 1882 1209
rect 1916 1175 1928 1209
rect 1870 1137 1928 1175
rect 1870 1103 1882 1137
rect 1916 1103 1928 1137
rect 1870 1065 1928 1103
rect 1870 1031 1882 1065
rect 1916 1031 1928 1065
rect 1870 993 1928 1031
rect 1870 959 1882 993
rect 1916 959 1928 993
rect 1870 921 1928 959
rect 1870 887 1882 921
rect 1916 887 1928 921
rect 1870 849 1928 887
rect 1870 815 1882 849
rect 1916 815 1928 849
rect 1870 777 1928 815
rect 1870 743 1882 777
rect 1916 743 1928 777
rect 1870 705 1928 743
rect 1870 671 1882 705
rect 1916 671 1928 705
rect 264 599 276 633
rect 310 599 322 633
rect 264 561 322 599
rect 264 527 276 561
rect 310 527 322 561
rect 264 489 322 527
rect 264 455 276 489
rect 310 455 322 489
rect 264 417 322 455
rect 264 383 276 417
rect 310 383 322 417
rect 264 322 322 383
rect 1870 633 1928 671
rect 1870 599 1882 633
rect 1916 599 1928 633
rect 1870 561 1928 599
rect 1870 527 1882 561
rect 1916 527 1928 561
rect 1870 489 1928 527
rect 1870 455 1882 489
rect 1916 455 1928 489
rect 1870 417 1928 455
rect 1870 383 1882 417
rect 1916 383 1928 417
rect 1870 322 1928 383
rect 264 310 1928 322
rect 264 276 276 310
rect 310 276 359 310
rect 393 276 431 310
rect 465 276 503 310
rect 537 276 575 310
rect 609 276 647 310
rect 681 276 719 310
rect 753 276 791 310
rect 825 276 863 310
rect 897 276 935 310
rect 969 276 1007 310
rect 1041 276 1079 310
rect 1113 276 1151 310
rect 1185 276 1223 310
rect 1257 276 1295 310
rect 1329 276 1367 310
rect 1401 276 1439 310
rect 1473 276 1511 310
rect 1545 276 1583 310
rect 1617 276 1655 310
rect 1689 276 1727 310
rect 1761 276 1799 310
rect 1833 276 1882 310
rect 1916 276 1928 310
rect 264 264 1928 276
rect 2096 3117 2154 3155
rect 2096 3083 2108 3117
rect 2142 3083 2154 3117
rect 2096 3045 2154 3083
rect 2096 3011 2108 3045
rect 2142 3011 2154 3045
rect 2096 2973 2154 3011
rect 2096 2939 2108 2973
rect 2142 2939 2154 2973
rect 2096 2901 2154 2939
rect 2096 2867 2108 2901
rect 2142 2867 2154 2901
rect 2096 2829 2154 2867
rect 2096 2795 2108 2829
rect 2142 2795 2154 2829
rect 2096 2757 2154 2795
rect 2096 2723 2108 2757
rect 2142 2723 2154 2757
rect 2096 2685 2154 2723
rect 2096 2651 2108 2685
rect 2142 2651 2154 2685
rect 2096 2613 2154 2651
rect 2096 2579 2108 2613
rect 2142 2579 2154 2613
rect 2096 2541 2154 2579
rect 2096 2507 2108 2541
rect 2142 2507 2154 2541
rect 2096 2469 2154 2507
rect 2096 2435 2108 2469
rect 2142 2435 2154 2469
rect 2096 2397 2154 2435
rect 2096 2363 2108 2397
rect 2142 2363 2154 2397
rect 2096 2325 2154 2363
rect 2096 2291 2108 2325
rect 2142 2291 2154 2325
rect 2096 2253 2154 2291
rect 2096 2219 2108 2253
rect 2142 2219 2154 2253
rect 2096 2181 2154 2219
rect 2096 2147 2108 2181
rect 2142 2147 2154 2181
rect 2096 2109 2154 2147
rect 2096 2075 2108 2109
rect 2142 2075 2154 2109
rect 2096 2037 2154 2075
rect 2096 2003 2108 2037
rect 2142 2003 2154 2037
rect 2096 1965 2154 2003
rect 2096 1931 2108 1965
rect 2142 1931 2154 1965
rect 2096 1893 2154 1931
rect 2096 1859 2108 1893
rect 2142 1859 2154 1893
rect 2096 1821 2154 1859
rect 2096 1787 2108 1821
rect 2142 1787 2154 1821
rect 2096 1749 2154 1787
rect 2096 1715 2108 1749
rect 2142 1715 2154 1749
rect 2096 1677 2154 1715
rect 2096 1643 2108 1677
rect 2142 1643 2154 1677
rect 2096 1605 2154 1643
rect 2096 1571 2108 1605
rect 2142 1571 2154 1605
rect 2096 1533 2154 1571
rect 2096 1499 2108 1533
rect 2142 1499 2154 1533
rect 2096 1461 2154 1499
rect 2096 1427 2108 1461
rect 2142 1427 2154 1461
rect 2096 1389 2154 1427
rect 2096 1355 2108 1389
rect 2142 1355 2154 1389
rect 2096 1317 2154 1355
rect 2096 1283 2108 1317
rect 2142 1283 2154 1317
rect 2096 1245 2154 1283
rect 2096 1211 2108 1245
rect 2142 1211 2154 1245
rect 2096 1173 2154 1211
rect 2096 1139 2108 1173
rect 2142 1139 2154 1173
rect 2096 1101 2154 1139
rect 2096 1067 2108 1101
rect 2142 1067 2154 1101
rect 2096 1029 2154 1067
rect 2096 995 2108 1029
rect 2142 995 2154 1029
rect 2096 957 2154 995
rect 2096 923 2108 957
rect 2142 923 2154 957
rect 2096 885 2154 923
rect 2096 851 2108 885
rect 2142 851 2154 885
rect 2096 813 2154 851
rect 2096 779 2108 813
rect 2142 779 2154 813
rect 2096 741 2154 779
rect 2096 707 2108 741
rect 2142 707 2154 741
rect 2096 669 2154 707
rect 2096 635 2108 669
rect 2142 635 2154 669
rect 2096 597 2154 635
rect 2096 563 2108 597
rect 2142 563 2154 597
rect 2096 525 2154 563
rect 2096 491 2108 525
rect 2142 491 2154 525
rect 2096 453 2154 491
rect 2096 419 2108 453
rect 2142 419 2154 453
rect 2096 381 2154 419
rect 2096 347 2108 381
rect 2142 347 2154 381
rect 2096 309 2154 347
rect 2096 275 2108 309
rect 2142 275 2154 309
rect 38 203 50 237
rect 84 203 96 237
rect 38 165 96 203
rect 38 131 50 165
rect 84 131 96 165
rect 38 96 96 131
rect 2096 237 2154 275
rect 2096 203 2108 237
rect 2142 203 2154 237
rect 2096 165 2154 203
rect 2096 131 2108 165
rect 2142 131 2154 165
rect 2096 96 2154 131
rect 38 84 2154 96
rect 38 50 50 84
rect 84 50 143 84
rect 177 50 215 84
rect 249 50 287 84
rect 321 50 359 84
rect 393 50 431 84
rect 465 50 503 84
rect 537 50 575 84
rect 609 50 647 84
rect 681 50 719 84
rect 753 50 791 84
rect 825 50 863 84
rect 897 50 935 84
rect 969 50 1007 84
rect 1041 50 1079 84
rect 1113 50 1151 84
rect 1185 50 1223 84
rect 1257 50 1295 84
rect 1329 50 1367 84
rect 1401 50 1439 84
rect 1473 50 1511 84
rect 1545 50 1583 84
rect 1617 50 1655 84
rect 1689 50 1727 84
rect 1761 50 1799 84
rect 1833 50 1871 84
rect 1905 50 1943 84
rect 1977 50 2015 84
rect 2049 50 2108 84
rect 2142 50 2154 84
rect 38 38 2154 50
<< properties >>
string GDS_END 9074670
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9004706
string path 7.850 12.350 7.850 76.950 46.950 76.950 46.950 7.850 3.350 7.850 
<< end >>
