magic
tech sky130A
magscale 1 2
timestamp 1679235063
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1383 203
rect 30 -17 64 21
<< locali >>
rect 17 289 337 323
rect 17 215 115 289
rect 161 215 269 255
rect 303 249 337 289
rect 1055 391 1105 493
rect 1223 391 1273 493
rect 1055 357 1273 391
rect 1223 331 1273 357
rect 303 215 379 249
rect 695 289 993 323
rect 695 265 729 289
rect 663 215 729 265
rect 763 215 887 255
rect 921 215 993 289
rect 1223 283 1384 331
rect 1322 181 1384 283
rect 1047 145 1384 181
rect 1047 55 1113 145
rect 1215 55 1281 145
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 27 391 77 493
rect 111 425 161 527
rect 195 391 245 493
rect 279 425 329 527
rect 363 459 581 493
rect 363 391 413 459
rect 531 427 581 459
rect 635 427 685 527
rect 719 459 937 493
rect 719 427 769 459
rect 27 357 413 391
rect 371 291 413 357
rect 447 393 497 425
rect 803 393 853 425
rect 447 283 524 393
rect 627 357 853 393
rect 887 357 937 459
rect 971 359 1021 527
rect 1139 433 1189 527
rect 1307 365 1357 527
rect 627 333 661 357
rect 591 299 661 333
rect 447 181 489 283
rect 591 249 629 299
rect 523 215 629 249
rect 1027 249 1092 323
rect 1027 215 1288 249
rect 591 181 629 215
rect 35 17 69 179
rect 103 95 153 181
rect 187 147 505 181
rect 187 129 254 147
rect 103 51 337 95
rect 371 17 405 111
rect 439 51 505 147
rect 591 145 945 181
rect 539 17 677 111
rect 711 51 777 145
rect 811 17 845 111
rect 879 51 945 145
rect 979 17 1013 179
rect 1147 17 1181 111
rect 1315 17 1349 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< obsm1 >>
rect 478 320 536 329
rect 1034 320 1092 329
rect 478 292 1092 320
rect 478 283 536 292
rect 1034 283 1092 292
<< labels >>
rlabel locali s 921 215 993 289 6 A1_N
port 1 nsew signal input
rlabel locali s 663 215 729 265 6 A1_N
port 1 nsew signal input
rlabel locali s 695 265 729 289 6 A1_N
port 1 nsew signal input
rlabel locali s 695 289 993 323 6 A1_N
port 1 nsew signal input
rlabel locali s 763 215 887 255 6 A2_N
port 2 nsew signal input
rlabel locali s 303 215 379 249 6 B1
port 3 nsew signal input
rlabel locali s 303 249 337 289 6 B1
port 3 nsew signal input
rlabel locali s 17 215 115 289 6 B1
port 3 nsew signal input
rlabel locali s 17 289 337 323 6 B1
port 3 nsew signal input
rlabel locali s 161 215 269 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 1383 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 1215 55 1281 145 6 X
port 9 nsew signal output
rlabel locali s 1047 55 1113 145 6 X
port 9 nsew signal output
rlabel locali s 1047 145 1384 181 6 X
port 9 nsew signal output
rlabel locali s 1322 181 1384 283 6 X
port 9 nsew signal output
rlabel locali s 1223 283 1384 331 6 X
port 9 nsew signal output
rlabel locali s 1223 331 1273 357 6 X
port 9 nsew signal output
rlabel locali s 1055 357 1273 391 6 X
port 9 nsew signal output
rlabel locali s 1223 391 1273 493 6 X
port 9 nsew signal output
rlabel locali s 1055 391 1105 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3926664
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3915260
<< end >>
